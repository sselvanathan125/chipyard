VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_io__analog_esd_pad
  CLASS PAD ;
  FOREIGN sky130_ef_io__analog_esd_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  PIN P_CORE
    PORT
      LAYER met3 ;
        RECT 24.720 0.000 49.720 82.350 ;
    END
  END P_CORE
  PIN VSSA
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
  END VSSA
  PIN VSSD
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
  END VSSD
  PIN AMUXBUS_B
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  PIN VDDIO_Q
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
  END VDDIO_Q
  PIN VDDIO
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
  END VDDIO
  PIN VSWITCH
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
  END VSWITCH
  PIN VSSIO
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.630 191.600 0.640 191.610 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.360 191.600 74.370 191.610 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
  END VSSIO
  PIN VDDA
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
  END VDDA
  PIN VCCD
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
  END VCCD
  PIN VCCHIB
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
  END VCCHIB
  PIN VSSIO_Q
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
  END VSSIO_Q
  PIN P_PAD
    PORT
      LAYER met5 ;
        RECT 7.050 105.120 67.890 165.945 ;
    END
  END P_PAD
  OBS
      LAYER li1 ;
        RECT 2.905 48.265 72.045 181.100 ;
      LAYER met1 ;
        RECT 4.250 46.255 70.440 48.855 ;
      LAYER met2 ;
        RECT 4.250 46.255 70.440 48.855 ;
      LAYER met3 ;
        RECT 0.455 82.750 74.250 173.315 ;
        RECT 0.455 14.905 24.320 82.750 ;
        RECT 50.120 14.905 74.250 82.750 ;
      LAYER met4 ;
        RECT 1.670 175.385 73.330 200.000 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 167.545 75.000 174.185 ;
        RECT 0.000 103.520 5.450 167.545 ;
        RECT 69.490 103.520 75.000 167.545 ;
        RECT 0.000 96.585 75.000 103.520 ;
        RECT 2.870 36.840 72.130 96.585 ;
        RECT 0.000 36.835 75.000 36.840 ;
        RECT 2.870 18.285 72.130 36.835 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_ef_io__analog_esd_pad

#--------EOF---------

MACRO sky130_ef_io__analog_noesd_pad
  CLASS PAD ;
  FOREIGN sky130_ef_io__analog_noesd_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  PIN P_CORE
    PORT
      LAYER met3 ;
        RECT 24.720 0.000 49.720 82.350 ;
    END
  END P_CORE
  PIN VSSA
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
  END VSSA
  PIN VSSD
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
  END VSSD
  PIN AMUXBUS_B
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  PIN VDDIO_Q
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
  END VDDIO_Q
  PIN VDDIO
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
  END VDDIO
  PIN VSWITCH
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
  END VSWITCH
  PIN VSSIO
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.630 191.600 0.640 191.610 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.360 191.600 74.370 191.610 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
  END VSSIO
  PIN VDDA
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
  END VDDA
  PIN VCCD
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
  END VCCD
  PIN VCCHIB
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
  END VCCHIB
  PIN VSSIO_Q
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
  END VSSIO_Q
  PIN P_PAD
    PORT
      LAYER met5 ;
        RECT 7.050 105.120 67.890 165.945 ;
    END
  END P_PAD
  OBS
      LAYER li1 ;
        RECT 2.905 48.265 72.045 181.100 ;
      LAYER met1 ;
        RECT 4.250 46.255 70.440 48.855 ;
      LAYER met2 ;
        RECT 4.250 46.255 70.440 48.855 ;
      LAYER met3 ;
        RECT 0.455 82.750 74.250 173.315 ;
        RECT 0.455 14.905 24.320 82.750 ;
        RECT 50.120 14.905 74.250 82.750 ;
      LAYER met4 ;
        RECT 1.670 175.385 73.330 200.000 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 167.545 75.000 174.185 ;
        RECT 0.000 103.520 5.450 167.545 ;
        RECT 69.490 103.520 75.000 167.545 ;
        RECT 0.000 96.585 75.000 103.520 ;
        RECT 2.870 36.840 72.130 96.585 ;
        RECT 0.000 36.835 75.000 36.840 ;
        RECT 2.870 18.285 72.130 36.835 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_ef_io__analog_noesd_pad

#--------EOF---------

MACRO sky130_ef_io__analog_pad
  CLASS PAD ;
  FOREIGN sky130_ef_io__analog_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  PIN P_CORE
    PORT
      LAYER met3 ;
        RECT 24.720 0.000 49.720 82.350 ;
    END
  END P_CORE
  PIN VSSA
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
  END VSSA
  PIN VSSD
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
  END VSSD
  PIN AMUXBUS_B
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  PIN VDDIO_Q
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
  END VDDIO_Q
  PIN VDDIO
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
  END VDDIO
  PIN VSWITCH
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
  END VSWITCH
  PIN VSSIO
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.630 191.600 0.640 191.610 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.360 191.600 74.370 191.610 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
  END VSSIO
  PIN VDDA
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
  END VDDA
  PIN VCCD
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
  END VCCD
  PIN VCCHIB
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
  END VCCHIB
  PIN VSSIO_Q
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
  END VSSIO_Q
  PIN P_PAD
    PORT
      LAYER met5 ;
        RECT 7.050 105.120 67.890 165.945 ;
    END
  END P_PAD
  OBS
      LAYER li1 ;
        RECT 2.905 48.265 72.045 181.100 ;
      LAYER met1 ;
        RECT 4.250 46.255 70.440 48.855 ;
      LAYER met2 ;
        RECT 4.250 46.255 70.440 48.855 ;
      LAYER met3 ;
        RECT 0.455 82.750 74.250 173.315 ;
        RECT 0.455 14.905 24.320 82.750 ;
        RECT 50.120 14.905 74.250 82.750 ;
      LAYER met4 ;
        RECT 1.670 175.385 73.330 200.000 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 167.545 75.000 174.185 ;
        RECT 0.000 103.520 5.450 167.545 ;
        RECT 69.490 103.520 75.000 167.545 ;
        RECT 0.000 96.585 75.000 103.520 ;
        RECT 2.870 36.840 72.130 96.585 ;
        RECT 0.000 36.835 75.000 36.840 ;
        RECT 2.870 18.285 72.130 36.835 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_ef_io__analog_pad

#--------EOF---------

MACRO sky130_ef_io__bare_pad
  CLASS BLOCK ;
  FOREIGN sky130_ef_io__bare_pad ;
  ORIGIN 2.700 2.700 ;
  SIZE 65.400 BY 75.400 ;
  PIN PAD
    PORT
      LAYER met4 ;
        RECT -2.700 70.000 62.700 72.700 ;
        RECT -2.700 0.000 0.000 70.000 ;
        RECT 60.000 0.000 62.700 70.000 ;
        RECT -2.700 -2.700 62.700 0.000 ;
      LAYER via4 ;
        RECT -2.580 71.400 62.580 72.580 ;
        RECT -2.580 -1.400 -1.400 71.400 ;
        RECT 61.400 -1.400 62.580 71.400 ;
        RECT -2.580 -2.580 62.580 -1.400 ;
      LAYER met5 ;
        RECT -2.700 -2.700 62.700 72.700 ;
    END
  END PAD
END sky130_ef_io__bare_pad

#--------EOF---------

MACRO sky130_ef_io__com_bus_slice_1um
  CLASS PAD SPACER ;
  FOREIGN sky130_ef_io__com_bus_slice_1um ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.800 1.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.000 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 1.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 1.000 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.000 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.000 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.000 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.000 92.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.000 22.400 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.000 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.750 1.000 197.965 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.000 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.000 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 0.000 173.75 1.000 197.965 ;
        RECT 0.000 66.900 1.000 67.600 ;
        RECT 0.000 61.050 1.000 61.650 ;
        RECT 0.000 55.100 1.000 55.800 ;
        RECT 0.000 49.610 1.000 50.790 ;
  END
END sky130_ef_io__com_bus_slice_1um

#--------EOF---------

MACRO sky130_ef_io__com_bus_slice_5um
  CLASS PAD SPACER ;
  FOREIGN sky130_ef_io__com_bus_slice_5um ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 5.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 5.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 5.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 5.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 5.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.800 5.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 5.000 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 5.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 5.000 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 5.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 5.000 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 5.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 5.000 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 5.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 5.000 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 5.000 92.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 5.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 5.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 5.000 22.400 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 5.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 5.000 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 5.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 5.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.750 5.000 197.965 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 5.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 5.000 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 5.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 5.000 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 0.000 173.75 5.000 197.965 ;
        RECT 0.000 66.900 5.000 67.600 ;
        RECT 0.000 61.050 5.000 61.650 ;
        RECT 0.000 55.100 5.000 55.800 ;
        RECT 0.000 49.610 5.000 50.790 ;
  END
END sky130_ef_io__com_bus_slice_5um

#--------EOF---------

MACRO sky130_ef_io__com_bus_slice_10um
  CLASS PAD SPACER ;
  FOREIGN sky130_ef_io__com_bus_slice_10um ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 10.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 10.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 10.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 10.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 10.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.800 10.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 10.000 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 10.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 10.000 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 10.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 10.000 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 10.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 10.000 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 10.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 10.000 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 10.000 92.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 10.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 10.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 10.000 22.400 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 10.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 10.000 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 10.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 10.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.750 10.000 197.965 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 10.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 10.000 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 10.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 10.000 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 0.000 173.75 10.000 197.965 ;
        RECT 0.000 66.900 10.000 67.600 ;
        RECT 0.000 61.050 10.000 61.650 ;
        RECT 0.000 55.100 10.000 55.800 ;
        RECT 0.000 49.610 10.000 50.790 ;
  END
END sky130_ef_io__com_bus_slice_10um

#--------EOF---------

MACRO sky130_ef_io__com_bus_slice_20um
  CLASS PAD SPACER ;
  FOREIGN sky130_ef_io__com_bus_slice_20um ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 20.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 20.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 20.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 20.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 20.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.800 20.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 20.000 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 20.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 20.000 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 20.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 20.000 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 20.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 20.000 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 20.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 20.000 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 20.000 92.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 20.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 20.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 20.000 22.400 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 20.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 20.000 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 20.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 20.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.750 20.000 197.965 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 20.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 20.000 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 20.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 20.000 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 0.000 173.75 20.000 197.965 ;
        RECT 0.000 66.900 20.000 67.600 ;
        RECT 0.000 61.050 20.000 61.650 ;
        RECT 0.000 55.100 20.000 55.800 ;
        RECT 0.000 49.610 20.000 50.790 ;
  END
END sky130_ef_io__com_bus_slice_20um

#--------EOF---------

MACRO sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
  CLASS PAD SPACER ;
  FOREIGN sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 20.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 20.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 20.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 20.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 20.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.800 20.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 20.000 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 20.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 20.000 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 20.000 33.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.990 17.880 19.000 33.200 ;
      LAYER via3 ;
        RECT 1.090 30.080 18.740 33.030 ;
        RECT 1.280 18.080 18.770 22.090 ;
      LAYER met4 ;
        RECT 0.000 29.850 20.000 33.300 ;
        RECT 0.000 17.750 20.000 22.400 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 20.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 20.000 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 20.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 20.000 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 20.000 92.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 20.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 20.000 22.300 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 20.000 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 20.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 20.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.750 20.000 197.965 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 20.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 20.000 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 20.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 20.000 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 0.000 173.750 20.000 197.965 ;
        RECT 0.000 49.610 20.000 50.790 ;
  END
END sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um

#--------EOF---------

MACRO sky130_ef_io__corner_pad
  CLASS ENDCAP TOPRIGHT ;
  FOREIGN sky130_ef_io__corner_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 204.000 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 57.125 22.910 60.105 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.125 0.000 56.105 26.910 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 52.365 20.935 55.345 ;
    END
    PORT
      LAYER met4 ;
        RECT 48.365 0.000 51.345 20.875 ;
    END
  END AMUXBUS_B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 51.735 23.155 60.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 40.835 1.335 44.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.735 19.575 52.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 40.735 1.335 44.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 55.645 21.550 56.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 60.405 23.175 60.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 36.840 0.000 40.085 1.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 47.735 0.000 56.735 27.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.405 0.000 56.735 27.175 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.645 0.000 52.825 21.555 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.735 0.000 40.185 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.735 0.000 48.065 23.575 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 19.035 1.470 22.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 18.935 1.470 22.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 15.035 0.000 18.285 1.255 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.935 0.000 18.385 1.255 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 35.985 1.385 39.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 35.885 1.385 39.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 31.985 0.000 35.235 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.885 0.000 35.335 1.270 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.185 1.480 72.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.085 1.480 72.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 64.185 0.000 68.435 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.085 0.000 68.535 1.270 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.135 2.350 11.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.035 2.350 11.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.135 0.000 7.385 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.035 0.000 7.485 1.270 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 74.035 2.645 98.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.885 1.525 28.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.785 1.525 28.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 74.035 2.645 99.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.885 0.000 24.335 1.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 70.035 0.000 94.985 1.855 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.035 0.000 95.000 1.855 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.785 0.000 24.435 1.270 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 12.985 3.785 17.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.885 3.785 17.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 8.985 0.000 13.435 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.885 0.000 13.535 1.270 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.935 1.600 34.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.835 1.600 34.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 179.785 1.435 204.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.935 0.000 30.385 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.835 0.000 30.485 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.785 0.000 200.000 1.270 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.685 1.475 50.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.585 1.475 50.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 41.685 0.000 46.135 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.585 0.000 46.235 1.270 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.335 1.625 66.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.235 1.625 66.685 ;
    END
    PORT
      LAYER met5 ;
        RECT 58.335 0.000 62.585 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.235 0.000 62.685 1.270 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 1.835 179.385 200.000 204.000 ;
        RECT 0.000 99.400 200.000 179.385 ;
        RECT 3.045 73.635 200.000 99.400 ;
        RECT 0.000 72.935 200.000 73.635 ;
        RECT 1.880 67.685 200.000 72.935 ;
        RECT 0.000 67.085 200.000 67.685 ;
        RECT 2.025 61.835 200.000 67.085 ;
        RECT 0.000 61.135 200.000 61.835 ;
        RECT 23.575 60.005 200.000 61.135 ;
        RECT 23.310 56.725 200.000 60.005 ;
        RECT 21.950 55.245 200.000 56.725 ;
        RECT 21.335 51.965 200.000 55.245 ;
        RECT 19.975 51.335 200.000 51.965 ;
        RECT 0.000 50.635 200.000 51.335 ;
        RECT 1.875 45.185 200.000 50.635 ;
        RECT 0.000 44.585 200.000 45.185 ;
        RECT 1.735 40.335 200.000 44.585 ;
        RECT 0.000 39.735 200.000 40.335 ;
        RECT 1.785 35.485 200.000 39.735 ;
        RECT 0.000 34.885 200.000 35.485 ;
        RECT 2.000 29.435 200.000 34.885 ;
        RECT 0.000 28.835 200.000 29.435 ;
        RECT 1.925 27.575 200.000 28.835 ;
        RECT 1.925 27.310 56.005 27.575 ;
        RECT 1.925 23.975 52.725 27.310 ;
        RECT 1.925 23.385 47.335 23.975 ;
        RECT 0.000 22.785 47.335 23.385 ;
        RECT 1.870 18.535 47.335 22.785 ;
        RECT 48.465 21.955 52.725 23.975 ;
        RECT 48.465 21.275 51.245 21.955 ;
        RECT 0.000 17.935 47.335 18.535 ;
        RECT 4.185 12.485 47.335 17.935 ;
        RECT 0.000 11.885 47.335 12.485 ;
        RECT 0.400 5.635 2.035 6.035 ;
        RECT 2.750 5.635 47.335 11.885 ;
        RECT 0.000 1.670 47.335 5.635 ;
        RECT 0.000 1.255 1.635 1.670 ;
        RECT 7.885 1.255 8.485 1.670 ;
        RECT 13.935 1.655 19.385 1.670 ;
        RECT 13.935 1.255 14.535 1.655 ;
        RECT 18.785 1.255 19.385 1.655 ;
        RECT 24.835 1.255 25.435 1.670 ;
        RECT 30.885 1.255 31.485 1.670 ;
        RECT 35.735 1.255 36.335 1.670 ;
        RECT 40.585 1.255 41.185 1.670 ;
        RECT 46.635 1.255 47.335 1.670 ;
        RECT 57.135 2.255 200.000 27.575 ;
        RECT 57.135 1.670 69.635 2.255 ;
        RECT 57.135 1.255 57.835 1.670 ;
        RECT 63.085 1.255 63.685 1.670 ;
        RECT 68.935 1.255 69.635 1.670 ;
        RECT 95.400 1.670 200.000 2.255 ;
        RECT 95.400 1.255 175.385 1.670 ;
      LAYER met5 ;
        RECT 0.000 100.585 200.000 204.000 ;
        RECT 4.245 72.435 200.000 100.585 ;
        RECT 3.080 68.185 200.000 72.435 ;
        RECT 3.225 62.335 200.000 68.185 ;
        RECT 24.755 50.135 200.000 62.335 ;
        RECT 3.075 44.085 200.000 50.135 ;
        RECT 2.935 40.835 200.000 44.085 ;
        RECT 2.985 35.985 200.000 40.835 ;
        RECT 3.200 28.755 200.000 35.985 ;
        RECT 3.200 28.335 46.135 28.755 ;
        RECT 3.125 22.285 46.135 28.335 ;
        RECT 3.070 19.035 46.135 22.285 ;
        RECT 5.385 11.385 46.135 19.035 ;
        RECT 1.600 4.535 2.135 6.135 ;
        RECT 3.950 4.535 46.135 11.385 ;
        RECT 0.000 2.870 46.135 4.535 ;
        RECT 58.335 3.455 200.000 28.755 ;
        RECT 58.335 2.870 68.435 3.455 ;
        RECT 0.000 0.000 0.535 2.870 ;
        RECT 15.035 2.855 18.285 2.870 ;
        RECT 96.585 0.000 200.000 3.455 ;
  END
END sky130_ef_io__corner_pad

#--------EOF---------

MACRO sky130_ef_io__disconnect_vccd_slice_5um
  CLASS PAD SPACER ;
  FOREIGN sky130_ef_io__disconnect_vccd_slice_5um ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 5.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 5.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 5.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 5.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 5.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.800 5.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 5.000 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 5.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 5.000 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 5.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 5.000 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 5.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 5.000 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 5.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 5.000 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 5.000 92.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 5.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 5.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 5.000 22.400 ;
    END
  END VDDIO
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 5.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 5.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.750 5.000 197.965 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 5.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 5.000 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 0.000 173.750 5.000 197.965 ;
        RECT 0.000 49.610 5.000 50.790 ;
  END
END sky130_ef_io__disconnect_vccd_slice_5um

#--------EOF---------

MACRO sky130_ef_io__disconnect_vdda_slice_5um
  CLASS PAD SPACER ;
  FOREIGN sky130_ef_io__disconnect_vdda_slice_5um ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 5.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 5.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 5.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 5.000 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 5.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 5.000 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 5.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 5.000 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 5.000 22.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 5.000 92.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 5.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 5.000 22.300 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 5.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 5.000 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 5.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 5.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.750 5.000 197.965 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 5.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 5.000 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 5.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 5.000 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 0.000 173.750 5.000 197.965 ;
  END
END sky130_ef_io__disconnect_vdda_slice_5um

#--------EOF---------

MACRO sky130_ef_io__gpiov2_pad
  CLASS PAD INOUT ;
  FOREIGN sky130_ef_io__gpiov2_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 36.440 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.760 51.090 80.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 52.145 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.465 46.330 80.000 49.310 ;
    END
  END AMUXBUS_B
  PIN ANALOG_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.430 -2.035 62.690 -0.730 ;
    END
  END ANALOG_EN
  PIN ANALOG_POL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.865 -2.035 46.195 34.770 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.750 -2.035 31.010 0.230 ;
    END
  END ANALOG_SEL
  PIN DM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.490 -2.035 28.750 2.035 ;
    END
  END DM[2]
  PIN DM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.835 -2.035 67.095 -0.840 ;
    END
  END DM[1]
  PIN DM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.855 -2.035 50.115 -1.490 ;
    END
  END DM[0]
  PIN ENABLE_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.460 -2.035 35.720 -0.485 ;
    END
  END ENABLE_H
  PIN ENABLE_INP_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.390 -2.035 38.650 1.055 ;
    END
  END ENABLE_INP_H
  PIN ENABLE_VDDA_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.755 -2.035 13.015 3.315 ;
    END
  END ENABLE_VDDA_H
  PIN ENABLE_VDDIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.580 -2.035 78.910 182.740 ;
    END
  END ENABLE_VDDIO
  PIN ENABLE_VSWITCH_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.310 -2.035 16.570 0.285 ;
    END
  END ENABLE_VSWITCH_H
  PIN HLD_H_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.815 -2.035 32.075 1.305 ;
    END
  END HLD_H_N
  PIN HLD_OVR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.600 -2.035 26.860 0.670 ;
    END
  END HLD_OVR
  PIN IB_MODE_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.420 -2.035 5.650 2.440 ;
    END
  END IB_MODE_SEL
  PIN IN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.240 -2.035 79.570 187.525 ;
    END
  END IN
  PIN IN_H
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.400 -2.035 1.020 176.450 ;
    END
  END IN_H
  PIN INP_DIS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.245 -2.035 45.505 3.055 ;
    END
  END INP_DIS
  PIN OE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.375 -2.035 3.605 2.440 ;
    END
  END OE_N
  PIN OUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.355 -2.035 22.615 4.390 ;
    END
  END OUT
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 11.200 102.525 73.800 164.975 ;
    END
  END PAD
  PIN PAD_A_ESD_0_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.280 -2.035 76.920 0.020 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.275 -2.035 68.925 0.235 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.820 -2.035 63.890 7.670 ;
    END
  END PAD_A_NOESD_H
  PIN SLOW
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.610 -2.035 77.870 -0.850 ;
    END
  END SLOW
  PIN TIE_HI_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.705 -2.035 78.905 -0.820 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.715 -2.035 79.915 175.835 ;
    END
  END TIE_LO_ESD
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 6.950 80.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 6.850 80.000 11.500 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 0.100 80.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 0.000 80.000 5.450 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.970 13.000 80.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.970 12.900 80.000 16.350 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 68.000 80.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 17.850 80.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 17.750 80.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 68.000 80.000 92.965 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 62.150 80.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 62.050 80.000 66.500 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 2.610 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 2.610 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 45.700 80.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 34.805 80.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 49.610 80.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.090 54.370 80.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.090 45.700 80.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 34.700 80.000 38.150 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 39.650 80.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 39.550 80.000 44.200 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 0.810 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.970 173.750 80.000 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 23.900 80.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 23.800 80.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 173.750 80.000 197.965 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 56.300 80.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 56.200 80.000 60.650 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 29.950 80.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 29.850 80.000 33.300 ;
    END
  END VSWITCH
  PIN VTRIP_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.130 -2.035 6.390 -0.485 ;
    END
  END VTRIP_SEL
  OBS
      LAYER nwell ;
        RECT -0.415 171.510 80.435 176.940 ;
        RECT -0.415 168.440 7.515 171.510 ;
        RECT 66.970 168.440 80.435 171.510 ;
        RECT -0.415 168.195 80.435 168.440 ;
        RECT -0.415 166.480 80.440 168.195 ;
        RECT -0.415 144.655 6.385 166.480 ;
        RECT 78.630 144.655 80.440 166.480 ;
        RECT -0.415 142.845 80.440 144.655 ;
      LAYER pwell ;
        RECT -0.290 138.650 80.290 142.530 ;
      LAYER nwell ;
        RECT 46.040 138.345 80.440 138.350 ;
        RECT -0.415 128.630 80.440 138.345 ;
      LAYER pwell ;
        RECT -0.215 127.280 40.245 128.320 ;
        RECT 66.910 127.280 80.290 128.320 ;
        RECT -0.215 123.100 80.290 127.280 ;
        RECT -0.215 101.515 5.735 123.100 ;
        RECT 77.865 101.515 80.290 123.100 ;
        RECT -0.215 99.930 80.290 101.515 ;
        RECT -0.215 94.220 5.215 99.930 ;
        RECT 39.385 98.785 80.290 99.930 ;
        RECT 52.880 97.485 80.290 98.785 ;
        RECT 76.770 95.950 80.290 97.485 ;
        RECT 39.385 94.220 80.290 95.950 ;
        RECT -0.215 93.940 80.290 94.220 ;
        RECT -0.215 93.225 45.840 93.940 ;
        RECT -0.215 92.920 46.590 93.225 ;
        RECT -0.215 90.900 9.300 92.920 ;
      LAYER nwell ;
        RECT 46.940 92.210 80.670 93.130 ;
        RECT 62.650 91.700 80.670 92.210 ;
        RECT -0.415 89.785 2.795 90.365 ;
        RECT -0.415 86.450 5.975 89.785 ;
        RECT -0.120 86.245 5.975 86.450 ;
        RECT -0.120 85.705 8.420 86.245 ;
        RECT -0.120 84.625 8.495 85.705 ;
        RECT -0.120 83.545 4.530 84.625 ;
        RECT 79.240 82.310 80.670 91.700 ;
        RECT 46.940 81.130 80.670 82.310 ;
        RECT -0.715 77.770 24.815 79.200 ;
        RECT -0.715 60.305 0.715 77.770 ;
        RECT 79.240 71.740 80.670 81.130 ;
        RECT 62.650 71.230 80.670 71.740 ;
        RECT 46.940 70.560 80.670 71.230 ;
        RECT 79.125 64.010 80.670 70.560 ;
        RECT 70.335 63.160 80.670 64.010 ;
        RECT -0.715 58.985 3.810 60.305 ;
        RECT -0.715 58.735 13.535 58.985 ;
        RECT -0.715 58.145 10.460 58.735 ;
        RECT -0.715 55.985 0.715 58.145 ;
        RECT -0.715 54.555 23.515 55.985 ;
        RECT 79.125 50.015 80.670 63.160 ;
        RECT 70.335 48.585 80.670 50.015 ;
        RECT 48.915 32.230 80.450 34.020 ;
        RECT 58.275 30.375 80.450 32.230 ;
        RECT 64.830 27.750 80.450 30.375 ;
        RECT 64.830 21.045 80.450 23.310 ;
        RECT 4.580 17.120 80.450 21.045 ;
        RECT -0.415 3.630 3.110 7.290 ;
        RECT 0.000 -2.035 61.490 1.465 ;
        RECT 64.030 -0.145 65.390 2.135 ;
      LAYER pwell ;
        RECT 64.245 -1.915 66.205 -0.905 ;
        RECT 66.610 -1.915 68.210 -0.655 ;
      LAYER li1 ;
        RECT 0.000 176.610 80.000 197.670 ;
        RECT -0.085 168.055 80.105 176.610 ;
        RECT -0.115 143.180 80.105 168.055 ;
        RECT -0.115 143.120 80.000 143.180 ;
        RECT 0.000 142.400 80.000 143.120 ;
        RECT -0.160 138.780 80.160 142.400 ;
        RECT 0.000 138.115 80.000 138.780 ;
        RECT -0.115 138.020 80.000 138.115 ;
        RECT -0.115 129.240 80.085 138.020 ;
        RECT -0.085 128.960 80.085 129.240 ;
        RECT 0.000 128.190 80.000 128.960 ;
        RECT -0.085 128.185 80.160 128.190 ;
        RECT -0.115 94.070 80.160 128.185 ;
        RECT -0.115 93.860 80.000 94.070 ;
        RECT -0.085 92.545 80.000 93.860 ;
        RECT -0.085 91.030 80.085 92.545 ;
        RECT 0.000 90.035 80.085 91.030 ;
        RECT -0.085 86.780 80.085 90.035 ;
        RECT 0.000 78.570 80.085 86.780 ;
        RECT -0.085 55.185 80.085 78.570 ;
        RECT 0.000 49.215 80.085 55.185 ;
        RECT 0.000 33.690 80.000 49.215 ;
        RECT 0.000 28.080 80.120 33.690 ;
        RECT 0.000 22.980 80.000 28.080 ;
        RECT 0.000 17.450 80.120 22.980 ;
        RECT 0.000 6.960 80.000 17.450 ;
        RECT -0.085 3.960 80.000 6.960 ;
        RECT 0.000 0.000 80.000 3.960 ;
        RECT 0.705 -0.100 0.875 0.000 ;
        RECT 0.705 -0.520 1.625 -0.100 ;
        RECT 2.090 -0.485 2.420 0.000 ;
        RECT 0.705 -1.500 0.875 -0.830 ;
        RECT 1.485 -0.860 1.655 -0.830 ;
        RECT 1.485 -1.390 1.660 -0.860 ;
        RECT 2.590 -1.345 2.760 0.000 ;
        RECT 3.470 -1.195 3.640 0.000 ;
        RECT 3.830 -0.080 4.160 0.000 ;
        RECT 4.350 -1.345 4.520 0.000 ;
        RECT 5.230 -1.195 5.400 0.000 ;
        RECT 6.110 -1.345 6.280 0.000 ;
        RECT 6.730 -1.345 6.900 0.000 ;
        RECT 7.610 -1.205 7.780 0.000 ;
        RECT 8.490 -1.345 8.660 0.000 ;
        RECT 9.370 -1.205 9.540 0.000 ;
        RECT 10.250 -1.345 10.420 0.000 ;
        RECT 10.615 -0.055 10.945 0.000 ;
        RECT 11.130 -1.205 11.300 0.000 ;
        RECT 11.750 -1.345 11.920 0.000 ;
        RECT 12.630 -1.205 12.800 0.000 ;
        RECT 13.510 -1.345 13.680 0.000 ;
        RECT 14.390 -1.205 14.560 0.000 ;
        RECT 15.270 -1.345 15.440 0.000 ;
        RECT 16.150 -1.205 16.320 0.000 ;
        RECT 17.030 -1.345 17.200 0.000 ;
        RECT 17.910 -1.205 18.080 0.000 ;
        RECT 18.790 -1.345 18.960 0.000 ;
        RECT 19.670 -1.205 19.840 0.000 ;
        RECT 20.550 -1.345 20.720 0.000 ;
        RECT 21.430 -1.205 21.600 0.000 ;
        RECT 22.310 -1.345 22.480 0.000 ;
        RECT 23.190 -1.205 23.360 0.000 ;
        RECT 24.070 -1.345 24.240 0.000 ;
        RECT 24.950 -1.205 25.120 0.000 ;
        RECT 25.830 -1.345 26.000 0.000 ;
        RECT 26.710 -1.205 26.880 0.000 ;
        RECT 27.590 -1.345 27.760 0.000 ;
        RECT 28.470 -1.205 28.640 0.000 ;
        RECT 29.350 -1.345 29.520 0.000 ;
        RECT 29.965 -0.050 30.495 0.000 ;
        RECT 29.970 -1.205 30.140 -0.050 ;
        RECT 30.850 -1.345 31.020 0.000 ;
        RECT 31.470 -1.345 31.640 0.000 ;
        RECT 32.350 -1.205 32.520 0.000 ;
        RECT 33.230 -1.345 33.400 0.000 ;
        RECT 34.110 -0.265 34.285 0.000 ;
        RECT 34.110 -1.205 34.280 -0.265 ;
        RECT 37.990 -1.345 38.160 0.000 ;
        RECT 38.870 -1.205 39.040 0.000 ;
        RECT 39.750 -1.345 39.920 0.000 ;
        RECT 40.630 -1.205 40.800 0.000 ;
        RECT 41.250 -1.345 41.420 0.000 ;
        RECT 42.130 -1.195 42.300 0.000 ;
        RECT 43.010 -1.345 43.180 0.000 ;
        RECT 45.290 -0.410 45.460 0.000 ;
        RECT 45.110 -0.580 45.640 -0.410 ;
        RECT 45.290 -1.205 45.460 -0.580 ;
        RECT 46.170 -1.345 46.340 0.000 ;
        RECT 47.050 -1.195 47.220 0.000 ;
        RECT 47.930 -1.345 48.100 0.000 ;
        RECT 48.495 -1.345 48.665 0.000 ;
        RECT 49.375 -1.205 49.545 0.000 ;
        RECT 50.255 -1.345 50.425 0.000 ;
        RECT 51.135 -1.205 51.305 0.000 ;
        RECT 52.015 -1.345 52.185 0.000 ;
        RECT 52.640 -1.205 52.810 0.000 ;
        RECT 53.520 -1.345 53.690 0.000 ;
        RECT 54.400 -1.205 54.570 0.000 ;
        RECT 54.750 -0.215 55.080 0.000 ;
        RECT 55.280 -1.345 55.450 0.000 ;
        RECT 55.830 -1.345 56.000 0.000 ;
        RECT 56.710 -1.205 56.880 0.000 ;
        RECT 57.590 -1.345 57.760 0.000 ;
        RECT 58.470 -1.205 58.640 0.000 ;
        RECT 59.020 -1.345 59.190 0.000 ;
        RECT 59.900 -1.205 60.070 0.000 ;
        RECT 60.780 -1.345 60.950 0.000 ;
        RECT 68.290 -0.095 70.005 0.000 ;
        RECT 72.315 -0.095 74.335 0.000 ;
        RECT 66.380 -0.575 67.270 -0.405 ;
        RECT 67.550 -0.575 68.220 -0.405 ;
        RECT 66.380 -0.795 66.910 -0.785 ;
        RECT 66.380 -0.955 66.965 -0.795 ;
        RECT 1.485 -1.500 1.655 -1.390 ;
        RECT 2.550 -1.705 60.990 -1.535 ;
        RECT 64.375 -1.785 66.075 -1.035 ;
        RECT 66.795 -1.805 66.965 -0.955 ;
        RECT 67.325 -1.805 67.495 -0.795 ;
        RECT 67.855 -0.815 68.025 -0.795 ;
        RECT 67.855 -0.985 68.385 -0.815 ;
        RECT 67.855 -1.805 68.025 -0.985 ;
      LAYER met1 ;
        RECT 0.000 178.940 80.000 197.965 ;
        RECT 0.000 176.865 80.020 178.940 ;
        RECT 0.000 168.055 80.000 176.865 ;
        RECT -0.115 129.240 80.145 168.055 ;
        RECT 0.000 128.185 80.000 129.240 ;
        RECT -0.115 93.860 80.145 128.185 ;
        RECT 0.000 92.545 80.000 93.860 ;
        RECT 0.000 89.445 80.060 92.545 ;
        RECT -0.145 87.715 80.060 89.445 ;
        RECT 0.000 78.600 80.060 87.715 ;
        RECT -0.115 70.895 80.060 78.600 ;
        POLYGON 80.060 70.950 80.115 70.895 80.060 70.895 ;
        RECT -0.115 55.155 80.115 70.895 ;
        RECT 0.000 49.185 80.115 55.155 ;
        RECT 0.000 33.690 80.000 49.185 ;
        RECT 0.000 28.085 80.115 33.690 ;
        RECT 0.000 22.980 80.000 28.085 ;
        RECT 0.000 17.450 80.115 22.980 ;
        RECT 0.000 0.000 80.000 17.450 ;
        RECT 0.260 -0.130 0.520 0.000 ;
        POLYGON 1.045 -0.100 1.045 -0.130 1.015 -0.130 ;
        RECT 1.045 -0.130 1.275 0.000 ;
        POLYGON 1.015 -0.130 1.015 -0.240 0.905 -0.240 ;
        RECT 1.015 -0.200 1.275 -0.130 ;
        RECT 1.015 -0.240 1.235 -0.200 ;
        POLYGON 1.235 -0.200 1.275 -0.200 1.235 -0.240 ;
        POLYGON 0.905 -0.240 0.905 -0.470 0.675 -0.470 ;
        RECT 0.675 -1.465 0.905 -0.470 ;
        POLYGON 0.905 -0.240 1.235 -0.240 0.905 -0.570 ;
        RECT 1.460 -0.610 1.690 0.000 ;
        POLYGON 1.690 -0.235 2.065 -0.610 1.690 -0.610 ;
        RECT 2.140 -0.255 2.370 0.000 ;
        RECT 3.880 -0.080 30.555 0.000 ;
        POLYGON 33.830 0.000 33.910 0.000 33.910 -0.080 ;
        RECT 33.910 -0.080 34.315 0.000 ;
        POLYGON 22.755 -0.080 22.760 -0.080 22.760 -0.085 ;
        RECT 22.760 -0.085 23.425 -0.080 ;
        POLYGON 2.370 -0.085 2.540 -0.255 2.370 -0.255 ;
        POLYGON 22.760 -0.085 22.785 -0.085 22.785 -0.110 ;
        RECT 22.785 -0.110 23.425 -0.085 ;
        POLYGON 23.425 -0.080 23.455 -0.080 23.425 -0.110 ;
        POLYGON 33.910 -0.080 33.940 -0.080 33.940 -0.110 ;
        RECT 33.940 -0.110 34.315 -0.080 ;
        POLYGON 35.570 0.000 35.655 0.000 35.655 -0.085 ;
        RECT 35.655 -0.085 42.895 0.000 ;
        POLYGON 42.895 0.000 42.980 0.000 42.895 -0.085 ;
        POLYGON 43.390 0.000 43.390 -0.085 43.305 -0.085 ;
        RECT 43.390 -0.085 47.720 0.000 ;
        POLYGON 33.940 -0.110 34.085 -0.110 34.085 -0.255 ;
        RECT 2.140 -0.485 18.040 -0.255 ;
        POLYGON 17.370 -0.485 17.400 -0.485 17.400 -0.515 ;
        RECT 17.400 -0.515 18.040 -0.485 ;
        RECT 21.550 -0.540 29.630 -0.280 ;
        RECT 29.770 -0.535 32.915 -0.275 ;
        RECT 34.085 -0.325 34.315 -0.110 ;
        POLYGON 43.305 -0.085 43.305 -0.225 43.165 -0.225 ;
        RECT 43.305 -0.190 47.720 -0.085 ;
        RECT 43.305 -0.225 43.370 -0.190 ;
        RECT 35.460 -0.485 38.120 -0.225 ;
        POLYGON 43.165 -0.225 43.165 -0.350 43.040 -0.350 ;
        RECT 43.165 -0.350 43.370 -0.225 ;
        POLYGON 43.370 -0.190 43.530 -0.190 43.370 -0.350 ;
        POLYGON 47.580 -0.190 47.680 -0.190 47.680 -0.290 ;
        RECT 47.680 -0.290 47.720 -0.190 ;
        POLYGON 47.720 0.000 48.010 -0.290 47.720 -0.290 ;
        POLYGON 54.810 -0.120 54.810 -0.290 54.640 -0.290 ;
        RECT 54.810 -0.290 55.040 0.000 ;
        RECT 56.680 -0.145 56.910 0.000 ;
        POLYGON 47.680 -0.290 47.740 -0.290 47.740 -0.350 ;
        RECT 47.740 -0.350 55.040 -0.290 ;
        RECT 39.390 -0.610 43.110 -0.350 ;
        POLYGON 43.110 -0.350 43.370 -0.350 43.110 -0.610 ;
        RECT 45.040 -0.610 47.515 -0.350 ;
        POLYGON 47.740 -0.350 47.910 -0.350 47.910 -0.520 ;
        RECT 47.910 -0.520 55.040 -0.350 ;
        RECT 1.460 -0.750 2.065 -0.610 ;
        POLYGON 2.065 -0.610 2.205 -0.750 2.065 -0.750 ;
        RECT 62.430 -0.730 62.690 -0.120 ;
        RECT 63.680 -0.595 64.880 0.000 ;
        POLYGON 65.530 0.000 65.635 0.000 65.635 -0.105 ;
        RECT 1.460 -1.765 61.195 -0.750 ;
        RECT 65.635 -0.845 65.775 0.000 ;
        POLYGON 66.830 -0.080 66.830 -0.375 66.535 -0.375 ;
        RECT 66.830 -0.375 67.095 0.000 ;
        RECT 66.320 -0.605 67.095 -0.375 ;
        RECT 67.355 -0.375 67.495 0.000 ;
        POLYGON 68.000 0.000 68.080 0.000 68.080 -0.080 ;
        RECT 68.080 -0.080 68.215 0.000 ;
        POLYGON 68.215 0.000 68.295 -0.080 68.215 -0.080 ;
        POLYGON 68.080 -0.080 68.215 -0.080 68.215 -0.215 ;
        RECT 68.215 -0.215 68.295 -0.080 ;
        POLYGON 67.495 -0.215 67.655 -0.375 67.495 -0.375 ;
        POLYGON 68.215 -0.215 68.295 -0.215 68.295 -0.295 ;
        POLYGON 68.295 -0.080 68.510 -0.295 68.295 -0.295 ;
        POLYGON 68.295 -0.295 68.370 -0.295 68.370 -0.370 ;
        RECT 67.355 -0.605 68.155 -0.375 ;
        POLYGON 68.370 -0.605 68.370 -0.705 68.270 -0.705 ;
        RECT 68.370 -0.705 68.510 -0.295 ;
        POLYGON 65.775 -0.705 65.915 -0.845 65.775 -0.845 ;
        POLYGON 68.270 -0.705 68.270 -0.755 68.220 -0.755 ;
        RECT 68.270 -0.755 68.510 -0.705 ;
        POLYGON 66.320 -0.755 66.320 -0.845 66.230 -0.845 ;
        RECT 66.320 -0.845 66.970 -0.755 ;
        POLYGON 68.220 -0.755 68.220 -0.785 68.190 -0.785 ;
        RECT 68.220 -0.785 68.510 -0.755 ;
        RECT 65.635 -0.985 66.970 -0.845 ;
        RECT 67.795 -1.015 68.510 -0.785 ;
        POLYGON 79.110 -0.915 79.110 -1.015 79.010 -1.015 ;
        RECT 79.110 -1.015 79.370 -0.835 ;
        POLYGON 79.010 -1.015 79.010 -1.125 78.900 -1.125 ;
        RECT 79.010 -1.125 79.370 -1.015 ;
        RECT 64.375 -1.775 67.525 -1.125 ;
        POLYGON 78.900 -1.125 78.900 -1.195 78.830 -1.195 ;
        RECT 78.900 -1.195 79.370 -1.125 ;
        RECT 75.255 -1.475 79.370 -1.195 ;
      LAYER met2 ;
        RECT 0.210 176.115 79.915 197.965 ;
        RECT 0.210 4.670 79.435 176.115 ;
        RECT 0.210 3.595 22.075 4.670 ;
        RECT 0.210 2.720 12.475 3.595 ;
        RECT 0.210 0.000 3.095 2.720 ;
        RECT 3.885 0.000 5.140 2.720 ;
        RECT 5.930 0.000 12.475 2.720 ;
        RECT 13.295 0.565 22.075 3.595 ;
        RECT 13.295 0.000 16.030 0.565 ;
        RECT 16.850 0.000 22.075 0.565 ;
        RECT 22.895 3.335 79.435 4.670 ;
        RECT 22.895 2.315 44.965 3.335 ;
        RECT 22.895 0.950 28.210 2.315 ;
        RECT 22.895 0.150 26.320 0.950 ;
        RECT 22.785 0.000 26.320 0.150 ;
        RECT 27.140 0.000 28.210 0.950 ;
        RECT 29.030 1.585 44.965 2.315 ;
        RECT 29.030 0.510 31.535 1.585 ;
        RECT 29.030 0.000 30.470 0.510 ;
        RECT 31.290 0.000 31.535 0.510 ;
        RECT 32.355 1.335 44.965 1.585 ;
        RECT 32.355 0.720 38.110 1.335 ;
        RECT 32.355 0.000 38.120 0.720 ;
        RECT 38.930 0.000 44.965 1.335 ;
        RECT 45.785 0.515 79.435 3.335 ;
        RECT 45.785 0.000 67.995 0.515 ;
        RECT 69.205 0.300 79.435 0.515 ;
        RECT 69.205 0.000 76.000 0.300 ;
        RECT 77.200 0.020 79.435 0.300 ;
        RECT 76.920 0.000 79.435 0.020 ;
        RECT 0.260 -1.065 0.520 0.000 ;
        RECT 1.080 -0.340 1.380 0.000 ;
        POLYGON 1.380 0.000 1.720 -0.340 1.380 -0.340 ;
        POLYGON 0.260 -1.065 0.520 -1.065 0.520 -1.325 ;
        POLYGON 0.520 -0.955 0.680 -1.115 0.520 -1.115 ;
        RECT 1.080 -1.110 1.720 -0.340 ;
        RECT 0.520 -1.325 0.680 -1.115 ;
        POLYGON 0.520 -1.325 0.670 -1.325 0.670 -1.475 ;
        RECT 0.670 -1.475 0.680 -1.325 ;
        POLYGON 0.680 -1.115 1.040 -1.475 0.680 -1.475 ;
        POLYGON 0.670 -1.475 0.930 -1.475 0.930 -1.735 ;
        RECT 0.930 -1.735 2.160 -1.475 ;
        RECT 2.365 -1.735 3.005 0.000 ;
        POLYGON 6.615 0.000 6.615 -0.020 6.595 -0.020 ;
        RECT 6.615 -0.020 6.965 0.000 ;
        POLYGON 6.965 0.000 6.985 0.000 6.965 -0.020 ;
        POLYGON 6.595 -0.020 6.595 -0.390 6.225 -0.390 ;
        POLYGON 6.595 -0.020 6.965 -0.020 6.595 -0.390 ;
        POLYGON 17.600 -0.080 17.600 -0.255 17.425 -0.255 ;
        RECT 17.600 -0.255 17.860 0.000 ;
        POLYGON 17.860 -0.080 18.035 -0.255 17.860 -0.255 ;
        POLYGON 6.225 -0.390 6.225 -0.485 6.130 -0.485 ;
        RECT 6.225 -0.485 6.500 -0.390 ;
        POLYGON 6.500 -0.390 6.595 -0.390 6.500 -0.485 ;
        POLYGON 6.390 -0.485 6.500 -0.485 6.390 -0.595 ;
        RECT 17.400 -0.515 18.040 -0.255 ;
        RECT 6.895 -1.765 10.715 -0.755 ;
        RECT 19.235 -1.765 21.375 0.000 ;
        POLYGON 21.775 -0.110 21.775 -0.280 21.605 -0.280 ;
        RECT 21.775 -0.280 22.035 0.000 ;
        RECT 22.785 -0.110 23.425 0.000 ;
        POLYGON 24.045 0.000 24.045 -0.110 23.935 -0.110 ;
        RECT 24.045 -0.110 26.265 0.000 ;
        POLYGON 23.935 -0.110 23.935 -0.125 23.920 -0.125 ;
        RECT 23.935 -0.125 26.265 -0.110 ;
        POLYGON 22.035 -0.125 22.190 -0.280 22.035 -0.280 ;
        POLYGON 23.920 -0.125 23.920 -0.150 23.895 -0.150 ;
        RECT 23.920 -0.150 26.265 -0.125 ;
        RECT 21.550 -0.540 22.190 -0.280 ;
        POLYGON 23.895 -0.150 23.895 -0.350 23.695 -0.350 ;
        RECT 23.895 -0.350 26.265 -0.150 ;
        POLYGON 23.695 -0.350 23.695 -0.540 23.505 -0.540 ;
        RECT 23.695 -0.540 26.265 -0.350 ;
        POLYGON 29.085 -0.185 29.085 -0.280 28.990 -0.280 ;
        RECT 29.085 -0.280 29.350 0.000 ;
        POLYGON 29.350 0.000 29.630 -0.280 29.350 -0.280 ;
        RECT 28.990 -0.540 29.630 -0.280 ;
        RECT 29.770 -0.535 30.410 0.000 ;
        POLYGON 32.355 -0.085 32.355 -0.165 32.275 -0.165 ;
        RECT 32.355 -0.165 32.615 0.000 ;
        RECT 32.275 -0.275 32.615 -0.165 ;
        POLYGON 32.615 -0.085 32.805 -0.275 32.615 -0.275 ;
        RECT 32.275 -0.535 32.915 -0.275 ;
        POLYGON 23.505 -0.540 23.505 -0.750 23.295 -0.750 ;
        RECT 23.505 -0.750 26.265 -0.540 ;
        RECT 22.995 -1.760 26.265 -0.750 ;
        RECT 33.400 -1.765 34.670 0.000 ;
        POLYGON 35.325 0.000 35.350 0.000 35.350 -0.025 ;
        RECT 35.350 -0.025 35.695 0.000 ;
        POLYGON 35.695 0.000 35.720 -0.025 35.695 -0.025 ;
        POLYGON 37.705 0.000 37.705 -0.025 37.680 -0.025 ;
        RECT 37.705 -0.025 38.120 0.000 ;
        POLYGON 35.350 -0.025 35.460 -0.025 35.460 -0.135 ;
        RECT 35.460 -0.225 35.720 -0.025 ;
        POLYGON 35.720 -0.025 35.920 -0.225 35.720 -0.225 ;
        POLYGON 37.680 -0.025 37.680 -0.225 37.480 -0.225 ;
        RECT 37.680 -0.225 38.120 -0.025 ;
        RECT 35.460 -0.485 36.100 -0.225 ;
        RECT 37.480 -0.485 38.120 -0.225 ;
        POLYGON 39.770 -0.005 39.770 -0.350 39.425 -0.350 ;
        RECT 39.770 -0.350 40.030 0.000 ;
        POLYGON 42.060 0.000 42.060 -0.310 41.750 -0.310 ;
        RECT 42.060 -0.310 42.120 0.000 ;
        POLYGON 42.120 0.000 42.430 0.000 42.120 -0.310 ;
        POLYGON 47.375 -0.180 47.375 -0.310 47.245 -0.310 ;
        RECT 47.375 -0.310 47.515 0.000 ;
        RECT 49.395 -0.165 50.165 0.000 ;
        POLYGON 35.720 -0.485 35.920 -0.485 35.720 -0.685 ;
        RECT 39.390 -0.610 40.030 -0.350 ;
        POLYGON 41.750 -0.310 41.750 -0.610 41.450 -0.610 ;
        POLYGON 41.450 -0.610 41.450 -0.680 41.380 -0.680 ;
        RECT 41.450 -0.680 41.750 -0.610 ;
        POLYGON 41.750 -0.310 42.120 -0.310 41.750 -0.680 ;
        POLYGON 47.245 -0.310 47.245 -0.350 47.205 -0.350 ;
        RECT 47.245 -0.350 47.515 -0.310 ;
        RECT 46.770 -0.610 47.515 -0.350 ;
        POLYGON 51.970 -0.330 51.970 -0.570 51.730 -0.570 ;
        RECT 51.970 -0.570 52.230 0.000 ;
        RECT 52.525 -0.040 54.155 0.000 ;
        POLYGON 52.525 -0.040 52.825 -0.040 52.825 -0.340 ;
        RECT 52.825 -0.340 54.155 -0.040 ;
        POLYGON 52.230 -0.340 52.460 -0.570 52.230 -0.570 ;
        POLYGON 41.380 -0.680 41.380 -0.685 41.375 -0.685 ;
        RECT 41.380 -0.685 41.530 -0.680 ;
        POLYGON 41.375 -0.685 41.375 -0.705 41.355 -0.705 ;
        RECT 41.375 -0.705 41.530 -0.685 ;
        POLYGON 38.650 -0.705 38.845 -0.900 38.650 -0.900 ;
        POLYGON 41.355 -0.705 41.355 -0.900 41.160 -0.900 ;
        RECT 41.355 -0.900 41.530 -0.705 ;
        POLYGON 41.530 -0.680 41.750 -0.680 41.530 -0.900 ;
        RECT 51.690 -0.850 52.460 -0.570 ;
        POLYGON 52.825 -0.340 53.335 -0.340 53.335 -0.850 ;
        RECT 53.335 -0.850 54.155 -0.340 ;
        POLYGON 53.335 -0.850 53.385 -0.850 53.385 -0.900 ;
        RECT 53.385 -0.900 54.155 -0.850 ;
        RECT 38.650 -1.160 41.270 -0.900 ;
        POLYGON 41.270 -0.900 41.530 -0.900 41.270 -1.160 ;
        POLYGON 53.385 -0.900 53.645 -0.900 53.645 -1.160 ;
        RECT 53.645 -0.985 54.155 -0.900 ;
        POLYGON 54.155 -0.185 54.955 -0.985 54.155 -0.985 ;
        RECT 62.430 -0.760 62.690 0.000 ;
        RECT 63.680 -0.595 64.385 0.000 ;
        POLYGON 76.920 0.000 77.330 0.000 76.920 -0.410 ;
        RECT 66.540 -0.840 67.360 -0.560 ;
        POLYGON 66.540 -0.840 66.685 -0.840 66.685 -0.985 ;
        RECT 66.685 -0.985 66.835 -0.840 ;
        RECT 53.645 -1.160 65.200 -0.985 ;
        POLYGON 66.685 -0.985 66.835 -0.985 66.835 -1.135 ;
        POLYGON 67.095 -0.840 67.360 -0.840 67.095 -1.105 ;
        RECT 77.390 -0.850 78.210 -0.570 ;
        POLYGON 78.710 -0.815 78.710 -0.820 78.705 -0.820 ;
        RECT 78.710 -0.820 78.910 0.000 ;
        POLYGON 77.410 -0.850 77.610 -0.850 77.610 -1.050 ;
        RECT 77.870 -1.050 77.980 -0.850 ;
        POLYGON 77.980 -0.850 78.180 -0.850 77.980 -1.050 ;
        RECT 78.905 -0.905 78.910 -0.820 ;
        POLYGON 78.905 -0.905 78.910 -0.905 78.905 -0.910 ;
        RECT 77.870 -1.105 77.925 -1.050 ;
        POLYGON 77.925 -1.050 77.980 -1.050 77.925 -1.105 ;
        RECT 77.870 -1.135 77.895 -1.105 ;
        POLYGON 77.895 -1.105 77.925 -1.105 77.895 -1.135 ;
        POLYGON 77.870 -1.135 77.895 -1.135 77.870 -1.160 ;
        POLYGON 38.650 -1.160 38.845 -1.160 38.650 -1.355 ;
        POLYGON 53.645 -1.160 53.695 -1.160 53.695 -1.210 ;
        RECT 53.695 -1.210 65.200 -1.160 ;
        RECT 49.590 -1.490 50.360 -1.210 ;
        POLYGON 49.590 -1.490 49.855 -1.490 49.855 -1.755 ;
        POLYGON 50.115 -1.490 50.360 -1.490 50.115 -1.735 ;
        POLYGON 53.695 -1.210 54.155 -1.210 54.155 -1.670 ;
        RECT 54.155 -1.670 65.200 -1.210 ;
        RECT 75.125 -1.475 75.895 -1.195 ;
        RECT 79.110 -1.475 79.370 0.000 ;
        POLYGON 54.155 -1.670 54.220 -1.670 54.220 -1.735 ;
        RECT 54.220 -1.735 65.200 -1.670 ;
        POLYGON 54.220 -1.735 54.240 -1.735 54.240 -1.755 ;
        RECT 54.240 -1.755 65.200 -1.735 ;
        POLYGON 54.240 -1.755 54.250 -1.755 54.250 -1.765 ;
        RECT 54.250 -1.765 65.200 -1.755 ;
        POLYGON 54.250 -1.765 54.270 -1.765 54.270 -1.785 ;
        RECT 54.270 -1.785 65.200 -1.765 ;
      LAYER met3 ;
        RECT 0.400 187.925 79.570 197.965 ;
        RECT 0.400 183.140 78.840 187.925 ;
        RECT 0.400 176.850 78.180 183.140 ;
        RECT 1.420 35.170 78.180 176.850 ;
        RECT 1.420 0.000 45.465 35.170 ;
        RECT 46.595 8.070 78.180 35.170 ;
        RECT 46.595 0.000 62.420 8.070 ;
        RECT 64.290 0.000 78.180 8.070 ;
        RECT 1.415 -1.090 2.205 -0.360 ;
        POLYGON 3.680 -1.125 3.680 -1.175 3.630 -1.175 ;
        RECT 3.680 -1.175 4.010 0.000 ;
        POLYGON 4.010 -0.775 4.410 -1.175 4.010 -1.175 ;
        RECT 3.630 -1.495 4.410 -1.175 ;
        RECT 6.455 -1.790 10.715 0.000 ;
        RECT 22.635 -1.785 27.635 0.000 ;
        RECT 49.415 -0.190 53.035 0.000 ;
        POLYGON 53.035 0.000 53.225 -0.190 53.035 -0.190 ;
        POLYGON 52.755 -0.190 53.110 -0.190 53.110 -0.545 ;
        RECT 53.110 -0.545 53.225 -0.190 ;
        POLYGON 53.225 -0.190 53.580 -0.545 53.225 -0.545 ;
        POLYGON 65.510 -0.310 65.510 -0.545 65.275 -0.545 ;
        RECT 65.510 -0.545 65.815 0.000 ;
        POLYGON 77.075 0.000 77.075 -0.415 76.660 -0.415 ;
        RECT 77.075 -0.415 77.110 0.000 ;
        POLYGON 77.110 0.000 77.525 0.000 77.110 -0.415 ;
        POLYGON 76.660 -0.415 76.660 -0.535 76.540 -0.535 ;
        RECT 51.685 -0.875 52.465 -0.545 ;
        POLYGON 53.110 -0.545 53.225 -0.545 53.225 -0.660 ;
        RECT 53.225 -0.660 54.320 -0.545 ;
        POLYGON 53.225 -0.660 53.430 -0.660 53.430 -0.865 ;
        RECT 53.430 -0.865 54.320 -0.660 ;
        POLYGON 55.510 -0.545 55.510 -0.865 55.190 -0.865 ;
        RECT 55.510 -0.865 56.785 -0.545 ;
        RECT 65.035 -0.865 65.815 -0.545 ;
        RECT 66.560 -0.865 67.340 -0.535 ;
        POLYGON 76.540 -0.535 76.540 -0.545 76.530 -0.545 ;
        RECT 76.540 -0.545 76.660 -0.535 ;
        RECT 75.120 -0.865 76.660 -0.545 ;
        POLYGON 76.660 -0.415 77.110 -0.415 76.660 -0.865 ;
        POLYGON 55.190 -0.865 55.190 -0.875 55.180 -0.875 ;
        RECT 55.190 -0.875 55.510 -0.865 ;
        POLYGON 55.180 -0.875 55.180 -0.995 55.060 -0.995 ;
        RECT 55.180 -0.995 55.510 -0.875 ;
        POLYGON 55.510 -0.865 55.640 -0.865 55.510 -0.995 ;
        RECT 77.410 -0.875 78.190 -0.545 ;
        POLYGON 55.060 -0.995 55.060 -1.185 54.870 -1.185 ;
        RECT 55.060 -1.185 55.205 -0.995 ;
        RECT 49.610 -1.300 55.205 -1.185 ;
        POLYGON 55.205 -0.995 55.510 -0.995 55.205 -1.300 ;
        RECT 49.610 -1.505 55.000 -1.300 ;
        POLYGON 55.000 -1.300 55.205 -1.300 55.000 -1.505 ;
        RECT 75.145 -1.500 75.925 -1.170 ;
        RECT 49.610 -1.515 50.340 -1.505 ;
        POLYGON 50.340 -1.505 50.350 -1.505 50.340 -1.515 ;
      LAYER met4 ;
        RECT 1.670 173.350 78.330 197.965 ;
        RECT 0.965 93.365 78.970 173.350 ;
        RECT 1.670 67.600 78.330 93.365 ;
        RECT 0.965 66.900 78.970 67.600 ;
        RECT 1.670 61.650 78.330 66.900 ;
        RECT 0.965 61.050 78.970 61.650 ;
        RECT 1.670 55.800 78.330 61.050 ;
        RECT 0.965 55.100 78.970 55.800 ;
        RECT 3.010 54.470 46.690 55.100 ;
        RECT 36.840 50.690 38.360 54.470 ;
        RECT 1.670 49.710 78.330 50.690 ;
        RECT 52.545 46.430 54.065 49.710 ;
        RECT 3.010 45.300 46.690 45.930 ;
        RECT 0.965 44.600 78.970 45.300 ;
        RECT 1.670 39.150 78.330 44.600 ;
        RECT 0.965 38.550 78.970 39.150 ;
        RECT 1.670 34.300 78.330 38.550 ;
        RECT 0.965 33.700 78.970 34.300 ;
        RECT 1.670 29.450 78.330 33.700 ;
        RECT 0.965 28.850 78.970 29.450 ;
        RECT 1.670 23.400 78.330 28.850 ;
        RECT 0.965 22.800 78.970 23.400 ;
        RECT 1.670 17.350 78.330 22.800 ;
        RECT 0.965 16.750 78.970 17.350 ;
        RECT 1.365 12.500 78.570 16.750 ;
        RECT 0.965 11.900 78.970 12.500 ;
        RECT 1.670 6.450 78.330 11.900 ;
        RECT 0.965 5.850 78.970 6.450 ;
        RECT 1.670 0.000 78.330 5.850 ;
        RECT 1.450 -0.870 52.440 -0.540 ;
        RECT 53.565 -0.870 56.760 -0.540 ;
        RECT 65.060 -0.870 67.315 -0.540 ;
        RECT 75.145 -0.870 78.165 -0.540 ;
        RECT 3.655 -1.500 75.900 -1.170 ;
      LAYER met5 ;
        RECT 0.000 166.575 80.000 197.965 ;
        RECT 0.000 100.925 9.600 166.575 ;
        RECT 75.400 100.925 80.000 166.575 ;
        RECT 0.000 94.550 80.000 100.925 ;
        RECT 2.870 16.250 77.130 94.550 ;
        RECT 2.565 13.000 77.370 16.250 ;
        RECT 2.870 0.100 77.130 13.000 ;
  END
END sky130_ef_io__gpiov2_pad

#--------EOF---------

MACRO sky130_ef_io__gpiov2_pad_wrapped
  CLASS PAD INOUT ;
  FOREIGN sky130_ef_io__gpiov2_pad_wrapped ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 210.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 64.090 36.440 67.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.760 64.090 80.000 67.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 59.330 52.145 62.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.465 59.330 80.000 62.310 ;
    END
  END AMUXBUS_B
  PIN ANALOG_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.705 0.000 50.985 2.400 ;
    END
  END ANALOG_EN
  PIN ANALOG_POL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.265 0.000 44.545 2.400 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.085 0.000 29.365 2.400 ;
    END
  END ANALOG_SEL
  PIN DM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.865 0.000 26.145 2.400 ;
    END
  END DM[2]
  PIN DM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.685 0.000 56.965 2.400 ;
    END
  END DM[1]
  PIN DM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.485 0.000 47.765 2.400 ;
    END
  END DM[0]
  PIN ENABLE_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.065 0.000 35.345 2.400 ;
    END
  END ENABLE_H
  PIN ENABLE_INP_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.285 0.000 38.565 2.400 ;
    END
  END ENABLE_INP_H
  PIN ENABLE_VDDA_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.445 0.000 13.725 2.400 ;
    END
  END ENABLE_VDDA_H
  PIN ENABLE_VDDIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.105 0.000 69.385 2.400 ;
    END
  END ENABLE_VDDIO
  PIN ENABLE_VSWITCH_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.665 0.000 16.945 2.400 ;
    END
  END ENABLE_VSWITCH_H
  PIN HLD_H_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.845 0.000 32.125 2.400 ;
    END
  END HLD_H_N
  PIN HLD_OVR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.645 0.000 22.925 2.400 ;
    END
  END HLD_OVR
  PIN IB_MODE_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.465 0.000 7.745 2.400 ;
    END
  END IB_MODE_SEL
  PIN IN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.085 0.000 75.365 2.400 ;
    END
  END IN
  PIN IN_H
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.485 0.000 1.765 2.400 ;
    END
  END IN_H
  PIN INP_DIS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.505 0.000 41.785 2.400 ;
    END
  END INP_DIS
  PIN OE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.245 0.000 4.525 2.400 ;
    END
  END OE_N
  PIN OUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.885 0.000 20.165 2.400 ;
    END
  END OUT
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 11.200 115.525 73.800 177.975 ;
    END
  END PAD
  PIN PAD_A_ESD_0_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.665 0.000 62.945 2.400 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.905 0.000 60.185 2.400 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.465 0.000 53.745 2.400 ;
    END
  END PAD_A_NOESD_H
  PIN SLOW
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.885 0.000 66.165 2.400 ;
    END
  END SLOW
  PIN TIE_HI_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.865 0.000 72.145 2.400 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.305 0.000 78.585 2.400 ;
    END
  END TIE_LO_ESD
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 19.950 1.270 24.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.850 1.270 24.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 19.950 80.000 24.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 19.850 80.000 24.500 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.100 1.270 18.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 13.000 1.270 18.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 13.100 80.000 18.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 13.000 80.000 18.450 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 26.000 0.965 29.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.900 0.965 29.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.970 26.000 80.000 29.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.970 25.900 80.000 29.350 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 81.000 1.270 105.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 30.850 1.270 35.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 30.750 1.270 35.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 81.000 1.270 105.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 81.000 80.000 105.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 30.850 80.000 35.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 30.750 80.000 35.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 81.000 80.000 105.965 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 75.150 1.270 79.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 75.050 1.270 79.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 75.150 80.000 79.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 75.050 80.000 79.500 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 58.700 1.270 67.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.805 1.270 51.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.700 2.610 59.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.610 1.270 63.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 67.370 2.610 67.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.700 1.270 51.150 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 58.700 80.000 67.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 47.805 80.000 51.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 62.610 80.000 63.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.090 67.370 80.000 67.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.090 58.700 80.000 59.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 47.700 80.000 51.150 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 52.650 1.270 57.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 52.550 1.270 57.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 52.650 80.000 57.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 52.550 80.000 57.200 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 186.750 1.270 210.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.900 1.270 41.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.800 1.270 41.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 186.750 80.000 210.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 36.900 80.000 41.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 36.800 80.000 41.450 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 69.300 1.270 73.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 69.200 1.270 73.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 69.300 80.000 73.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 69.200 80.000 73.650 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 42.950 1.270 46.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 42.850 1.270 46.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 42.950 80.000 46.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 42.850 80.000 46.300 ;
    END
  END VSWITCH
  PIN VTRIP_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.685 0.000 10.965 2.400 ;
    END
  END VTRIP_SEL
  OBS
      LAYER li1 ;
        RECT -0.160 11.195 80.160 210.670 ;
      LAYER met1 ;
        RECT -0.145 4.120 80.145 210.965 ;
      LAYER met2 ;
        RECT 0.210 2.680 79.915 210.965 ;
        RECT 0.210 2.400 1.205 2.680 ;
        RECT 2.045 2.400 3.965 2.680 ;
        RECT 4.805 2.400 7.185 2.680 ;
        RECT 8.025 2.400 10.405 2.680 ;
        RECT 11.245 2.400 13.165 2.680 ;
        RECT 14.005 2.400 16.385 2.680 ;
        RECT 17.225 2.400 19.605 2.680 ;
        RECT 20.445 2.400 22.365 2.680 ;
        RECT 23.205 2.400 25.585 2.680 ;
        RECT 26.425 2.400 28.805 2.680 ;
        RECT 29.645 2.400 31.565 2.680 ;
        RECT 32.405 2.400 34.785 2.680 ;
        RECT 35.625 2.400 38.005 2.680 ;
        RECT 38.845 2.400 41.225 2.680 ;
        RECT 42.065 2.400 43.985 2.680 ;
        RECT 44.825 2.400 47.205 2.680 ;
        RECT 48.045 2.400 50.425 2.680 ;
        RECT 51.265 2.400 53.185 2.680 ;
        RECT 54.025 2.400 56.405 2.680 ;
        RECT 57.245 2.400 59.625 2.680 ;
        RECT 60.465 2.400 62.385 2.680 ;
        RECT 63.225 2.400 65.605 2.680 ;
        RECT 66.445 2.400 68.825 2.680 ;
        RECT 69.665 2.400 71.585 2.680 ;
        RECT 72.425 2.400 74.805 2.680 ;
        RECT 75.645 2.400 78.025 2.680 ;
        RECT 78.865 2.400 79.915 2.680 ;
      LAYER met3 ;
        RECT 0.310 9.655 79.570 210.965 ;
      LAYER met4 ;
        RECT 1.670 186.350 78.330 210.965 ;
        RECT 0.965 106.365 78.970 186.350 ;
        RECT 1.670 80.600 78.330 106.365 ;
        RECT 0.965 79.900 78.970 80.600 ;
        RECT 1.670 74.650 78.330 79.900 ;
        RECT 0.965 74.050 78.970 74.650 ;
        RECT 1.670 68.800 78.330 74.050 ;
        RECT 0.965 68.100 78.970 68.800 ;
        RECT 3.010 67.470 46.690 68.100 ;
        RECT 36.840 63.690 38.360 67.470 ;
        RECT 1.670 62.710 78.330 63.690 ;
        RECT 52.545 59.430 54.065 62.710 ;
        RECT 3.010 58.300 46.690 58.930 ;
        RECT 0.965 57.600 78.970 58.300 ;
        RECT 1.670 52.150 78.330 57.600 ;
        RECT 0.965 51.550 78.970 52.150 ;
        RECT 1.670 47.300 78.330 51.550 ;
        RECT 0.965 46.700 78.970 47.300 ;
        RECT 1.670 42.450 78.330 46.700 ;
        RECT 0.965 41.850 78.970 42.450 ;
        RECT 1.670 36.400 78.330 41.850 ;
        RECT 0.965 35.800 78.970 36.400 ;
        RECT 1.670 30.350 78.330 35.800 ;
        RECT 0.965 29.750 78.970 30.350 ;
        RECT 1.365 25.500 78.570 29.750 ;
        RECT 0.965 24.900 78.970 25.500 ;
        RECT 1.670 19.450 78.330 24.900 ;
        RECT 0.965 18.850 78.970 19.450 ;
        RECT 1.670 12.600 78.330 18.850 ;
        RECT 0.965 11.500 78.970 12.600 ;
      LAYER met5 ;
        RECT 0.000 179.575 80.000 210.965 ;
        RECT 0.000 113.925 9.600 179.575 ;
        RECT 75.400 113.925 80.000 179.575 ;
        RECT 0.000 107.550 80.000 113.925 ;
        RECT 2.870 29.250 77.130 107.550 ;
        RECT 2.565 26.000 77.370 29.250 ;
        RECT 2.870 13.100 77.130 26.000 ;
  END
END sky130_ef_io__gpiov2_pad_wrapped

#--------EOF---------

MACRO sky130_ef_io__top_power_hvc
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__top_power_hvc ;
  ORIGIN 0.000 0.000 ;
  SIZE 169.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 169.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 169.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 97.390 -2.035 121.290 23.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.890 -2.035 95.890 9.295 ;
    END
  END DRN_HVC
  PIN P_CORE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 -2.035 71.395 13.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.390 -2.035 169.000 13.650 ;
    END
  END P_CORE
  PIN P_PAD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 54.050 103.085 114.890 163.910 ;
    END
  END P_PAD
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 47.495 -2.035 71.395 0.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.895 -2.035 83.895 0.690 ;
    END
  END SRC_BDY_HVC
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 125.885 45.700 169.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 125.885 34.800 169.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.885 49.610 169.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 169.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 169.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.885 34.700 169.000 38.150 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 47.240 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.800 47.715 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 47.240 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 47.715 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 121.205 13.000 169.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.205 12.900 169.000 16.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 47.715 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 47.715 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 125.885 29.950 169.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.885 29.850 169.000 33.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 47.715 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 47.715 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 125.885 62.150 169.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.885 62.050 169.000 66.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 47.715 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 47.715 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 125.885 0.100 169.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.885 0.000 169.000 5.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 47.715 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 47.715 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 125.885 68.000 169.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 125.885 17.850 169.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.205 17.750 169.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.885 68.000 169.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 47.715 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 47.715 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 47.715 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 47.715 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 125.885 6.950 169.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.885 6.850 169.000 11.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 47.715 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 47.715 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 128.245 173.750 169.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 168.360 189.565 168.370 189.575 ;
    END
    PORT
      LAYER met5 ;
        RECT 125.885 23.900 169.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.885 23.800 169.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 167.730 173.750 169.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 48.205 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.630 189.565 0.640 189.575 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 47.715 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 47.715 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 125.885 39.650 169.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.885 39.550 169.000 44.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 47.715 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 47.250 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 125.885 56.300 169.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.885 56.200 169.000 60.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 47.715 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 47.715 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER pwell ;
        RECT 50.495 -1.100 58.285 21.755 ;
      LAYER nwell ;
        RECT 58.860 -1.350 117.965 0.170 ;
      LAYER li1 ;
        RECT 47.610 0.000 119.855 197.660 ;
        RECT 47.610 -0.970 58.155 0.000 ;
        RECT 59.035 -0.115 60.045 0.000 ;
        RECT 116.730 -0.115 117.680 0.000 ;
        RECT 59.035 -1.065 117.680 -0.115 ;
      LAYER met1 ;
        RECT 47.185 0.000 119.915 197.690 ;
        RECT 50.625 -0.905 55.855 0.000 ;
        RECT 59.035 -0.115 60.350 0.000 ;
        POLYGON 60.350 0.000 60.465 -0.115 60.350 -0.115 ;
        POLYGON 116.540 0.000 116.540 -0.115 116.425 -0.115 ;
        RECT 116.540 -0.115 117.680 0.000 ;
        RECT 59.035 -1.065 117.680 -0.115 ;
      LAYER met2 ;
        RECT 47.265 23.905 121.290 193.040 ;
        RECT 47.265 0.300 97.110 23.905 ;
        RECT 71.675 0.000 97.110 0.300 ;
        RECT 72.895 -2.035 74.895 -0.115 ;
      LAYER met3 ;
        RECT 0.000 14.050 169.000 197.965 ;
        RECT 71.795 9.695 96.990 14.050 ;
        RECT 71.795 1.090 84.490 9.695 ;
        RECT 71.795 0.690 72.495 1.090 ;
        RECT 84.295 0.690 84.490 1.090 ;
        RECT 96.290 0.690 96.990 9.695 ;
      LAYER met4 ;
        RECT 48.605 173.350 127.845 197.965 ;
        RECT 47.240 93.365 128.245 173.350 ;
        RECT 48.115 67.600 125.485 93.365 ;
        RECT 47.240 66.900 128.245 67.600 ;
        RECT 48.115 61.650 125.485 66.900 ;
        RECT 47.240 61.050 128.245 61.650 ;
        RECT 48.115 55.800 125.485 61.050 ;
        RECT 47.240 55.100 128.245 55.800 ;
        RECT 47.640 49.710 125.485 50.690 ;
        RECT 47.240 44.600 128.245 45.300 ;
        RECT 47.650 39.150 125.485 44.600 ;
        RECT 47.240 38.550 128.245 39.150 ;
        RECT 48.115 34.300 125.485 38.550 ;
        RECT 47.240 33.700 128.245 34.300 ;
        RECT 48.115 29.450 125.485 33.700 ;
        RECT 47.240 28.850 128.245 29.450 ;
        RECT 48.115 23.400 125.485 28.850 ;
        RECT 47.240 22.800 128.245 23.400 ;
        RECT 48.115 17.350 120.805 22.800 ;
        RECT 47.240 16.750 128.245 17.350 ;
        RECT 48.115 12.500 120.805 16.750 ;
        RECT 47.240 11.900 128.245 12.500 ;
        RECT 48.115 6.450 125.485 11.900 ;
        RECT 47.240 5.850 128.245 6.450 ;
        RECT 48.115 0.000 125.485 5.850 ;
      LAYER met5 ;
        RECT 0.000 165.510 169.000 197.965 ;
        RECT 0.000 101.485 52.450 165.510 ;
        RECT 116.490 101.485 169.000 165.510 ;
        RECT 0.000 94.550 169.000 101.485 ;
        RECT 49.315 54.700 124.285 94.550 ;
        RECT 48.840 45.700 124.285 54.700 ;
        RECT 49.315 17.850 124.285 45.700 ;
        RECT 49.315 11.400 119.605 17.850 ;
        RECT 49.315 0.100 124.285 11.400 ;
  END
END sky130_ef_io__top_power_hvc

#--------EOF---------

MACRO sky130_ef_io__vccd_hvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vccd_hvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 50.390 -2.035 74.290 23.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 -2.035 48.890 9.295 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.495 -2.035 24.395 0.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895 -2.035 36.895 0.690 ;
    END
  END SRC_BDY_HVC
  PIN VCCD_PAD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 7.050 103.085 67.890 163.910 ;
    END
  END VCCD_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 6.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 6.865 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER pwell ;
        RECT 3.495 -1.100 11.285 21.755 ;
      LAYER nwell ;
        RECT 11.860 -1.350 70.965 0.170 ;
      LAYER li1 ;
        RECT 0.610 0.000 72.855 197.660 ;
        RECT 0.610 -0.970 11.155 0.000 ;
        RECT 12.035 -0.115 13.045 0.000 ;
        RECT 69.730 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met1 ;
        RECT 0.185 0.000 72.915 197.690 ;
        RECT 3.625 -0.905 8.855 0.000 ;
        RECT 12.035 -0.115 13.350 0.000 ;
        POLYGON 13.350 0.000 13.465 -0.115 13.350 -0.115 ;
        POLYGON 69.540 0.000 69.540 -0.115 69.425 -0.115 ;
        RECT 69.540 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met2 ;
        RECT 0.265 23.905 74.290 193.040 ;
        RECT 0.265 0.300 50.110 23.905 ;
        RECT 24.675 0.000 50.110 0.300 ;
        RECT 25.895 -2.035 27.895 -0.115 ;
      LAYER met3 ;
        RECT 0.240 9.695 74.290 197.965 ;
        RECT 0.240 7.265 37.490 9.695 ;
        RECT 24.795 1.090 37.490 7.265 ;
        RECT 24.795 0.690 25.495 1.090 ;
        RECT 37.295 0.690 37.490 1.090 ;
        RECT 49.290 7.265 74.290 9.695 ;
        RECT 49.290 0.690 49.990 7.265 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 165.510 75.000 197.965 ;
        RECT 0.000 101.485 5.450 165.510 ;
        RECT 69.490 101.485 75.000 165.510 ;
        RECT 0.000 94.550 75.000 101.485 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vccd_hvc_pad

#--------EOF---------

MACRO sky130_ef_io__vccd_lvc_clamped2_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vccd_lvc_clamped2_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN VCCD_PAD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 10.270 99.865 64.670 167.130 ;
    END
  END VCCD_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 6.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 6.865 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 76.470 197.930 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 75.000 197.805 ;
        RECT 16.655 -0.035 56.565 0.000 ;
        RECT 20.925 -0.815 56.565 -0.035 ;
        RECT 76.200 -0.815 85.935 75.350 ;
        RECT 20.925 -6.920 85.935 -0.815 ;
        RECT 20.925 -10.920 81.935 -6.920 ;
        POLYGON 81.935 -6.920 85.935 -6.920 81.935 -10.920 ;
      LAYER met2 ;
        RECT 0.000 44.200 75.000 197.930 ;
        RECT 76.200 46.560 85.935 197.930 ;
        RECT 0.000 44.165 86.140 44.200 ;
        RECT -10.975 39.550 86.140 44.165 ;
        RECT -10.975 39.515 75.000 39.550 ;
        RECT 0.000 0.000 75.000 39.515 ;
        RECT 76.200 23.390 85.935 37.800 ;
        RECT 0.500 -0.035 20.495 0.000 ;
        RECT 20.925 -0.035 53.535 0.000 ;
        RECT 54.095 -0.035 74.700 0.000 ;
      LAYER met3 ;
        RECT -10.975 39.515 -0.895 44.165 ;
        RECT 0.000 7.265 75.000 197.930 ;
        RECT 76.200 173.715 85.935 197.930 ;
        RECT 75.605 39.550 86.140 44.200 ;
        RECT 76.200 23.765 85.935 28.415 ;
        RECT 0.000 0.000 0.100 7.265 ;
        RECT 24.900 0.000 50.355 7.265 ;
        RECT 26.000 -0.035 36.880 0.000 ;
        RECT 38.380 -0.035 49.255 0.000 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 76.470 173.750 85.935 197.930 ;
        RECT 74.785 173.715 85.935 173.750 ;
        RECT 0.000 93.365 75.000 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.000 66.900 75.000 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.000 61.050 75.000 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.000 55.100 75.000 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.000 44.600 75.000 45.300 ;
        RECT -10.975 39.550 0.000 44.165 ;
        RECT -10.975 39.515 0.070 39.550 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 75.000 39.550 86.140 44.200 ;
        RECT 0.000 38.550 75.000 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.000 33.700 75.000 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.000 28.850 75.000 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 75.000 23.800 85.935 28.415 ;
        RECT 74.935 23.765 85.935 23.800 ;
        RECT 0.000 22.800 75.000 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.000 16.750 75.000 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.000 11.900 75.000 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.000 5.850 75.000 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 168.730 75.000 197.965 ;
        RECT 0.000 98.265 8.670 168.730 ;
        RECT 66.270 98.265 75.000 168.730 ;
        RECT 0.000 94.550 75.000 98.265 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vccd_lvc_clamped2_pad

#--------EOF---------

MACRO sky130_ef_io__vccd_lvc_clamped3_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vccd_lvc_clamped3_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VCCD_PAD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 10.270 99.865 64.670 167.130 ;
    END
  END VCCD_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 76.470 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  PIN VCCD1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER met3 ;
        RECT 0.500 -7.830 24.500 47.345 ;
    END
    PORT
      CLASS CORE ;
      LAYER met3 ;
        RECT 50.755 -7.710 74.700 84.430 ;
    END
  END VCCD1
  PIN VSSD1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER met3 ;
        RECT 25.950 -7.530 49.260 -2.510 ;
    END
  END VSSD1
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 75.000 197.805 ;
        RECT 16.655 -0.035 56.565 0.000 ;
        RECT 20.925 -0.780 56.565 -0.035 ;
        RECT 76.200 -0.780 85.935 75.385 ;
        RECT 20.925 -6.885 85.935 -0.780 ;
        RECT 20.925 -10.885 81.935 -6.885 ;
        POLYGON 81.935 -6.885 85.935 -6.885 81.935 -10.885 ;
      LAYER met2 ;
        RECT 0.490 0.000 75.000 197.965 ;
        RECT 76.200 23.425 85.935 197.965 ;
        RECT 0.490 -2.510 20.495 0.000 ;
        RECT 20.925 -0.035 53.535 0.000 ;
        POLYGON 20.495 -1.510 21.495 -2.510 20.495 -2.510 ;
        POLYGON 54.095 -1.510 54.095 -2.510 53.095 -2.510 ;
        RECT 54.095 -2.510 74.700 0.000 ;
        RECT 0.490 -2.560 74.700 -2.510 ;
        POLYGON 0.490 -2.560 5.490 -2.560 5.490 -7.560 ;
        RECT 5.490 -7.560 69.700 -2.560 ;
        POLYGON 69.700 -2.560 74.700 -2.560 69.700 -7.560 ;
      LAYER met3 ;
        RECT 0.490 84.830 75.000 197.965 ;
        RECT 76.200 173.750 85.935 197.965 ;
        RECT 0.490 47.745 50.355 84.830 ;
        RECT 0.490 -7.830 0.500 4.310 ;
        RECT 24.900 0.000 50.355 47.745 ;
        RECT 76.200 23.800 85.935 28.450 ;
        RECT 26.000 -0.035 36.880 0.000 ;
        RECT 38.380 -0.035 49.255 0.000 ;
      LAYER met4 ;
        RECT 1.605 173.350 73.825 197.965 ;
        RECT 76.470 173.750 85.935 197.965 ;
        RECT 0.965 93.365 75.000 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 75.000 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 75.000 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 75.000 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 75.000 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 75.000 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 75.000 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 75.000 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 75.000 23.800 85.935 28.450 ;
        RECT 0.965 22.800 75.000 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 75.000 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 75.000 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 75.000 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 168.730 75.000 197.965 ;
        RECT 0.000 98.265 8.670 168.730 ;
        RECT 66.270 98.265 75.000 168.730 ;
        RECT 0.000 94.550 75.000 98.265 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vccd_lvc_clamped3_pad

#--------EOF---------

MACRO sky130_ef_io__vccd_lvc_clamped_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vccd_lvc_clamped_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN VCCD_PAD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 10.270 99.865 64.670 167.130 ;
    END
  END VCCD_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 6.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 6.865 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 0.705 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 75.000 197.805 ;
        RECT 75.245 34.455 86.195 38.325 ;
        RECT 16.655 -0.035 56.565 0.000 ;
        RECT 20.495 -0.815 56.565 -0.035 ;
        RECT 76.200 -0.815 85.935 34.455 ;
        RECT 20.495 -1.015 85.935 -0.815 ;
        POLYGON 18.655 -1.015 18.655 -3.015 16.655 -3.015 ;
        RECT 18.655 -3.015 85.935 -1.015 ;
        RECT 16.655 -6.535 85.935 -3.015 ;
        RECT 16.655 -8.535 81.935 -6.535 ;
        POLYGON 16.655 -8.535 18.655 -8.535 18.655 -10.535 ;
        RECT 18.655 -10.535 81.935 -8.535 ;
        POLYGON 81.935 -6.535 85.935 -6.535 81.935 -10.535 ;
      LAYER met2 ;
        RECT 0.490 44.200 75.000 194.395 ;
        RECT 0.490 39.550 86.140 44.200 ;
        RECT 0.490 0.000 75.000 39.550 ;
        RECT 75.245 34.455 86.195 38.325 ;
        RECT 0.500 -0.035 20.495 0.000 ;
        RECT 20.925 -0.035 53.535 0.000 ;
        RECT 54.095 -0.035 74.700 0.000 ;
      LAYER met3 ;
        RECT 0.490 7.265 75.000 193.570 ;
        RECT 75.605 39.550 86.140 44.200 ;
        RECT 75.440 34.695 86.140 38.160 ;
        RECT 24.900 0.000 50.355 7.265 ;
        RECT 26.000 -0.035 36.880 0.000 ;
        RECT 38.380 -0.035 49.255 0.000 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 75.000 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 75.000 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 75.000 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 75.000 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 75.000 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 75.000 39.550 86.140 44.200 ;
        RECT 0.965 38.550 75.000 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 75.000 34.700 86.165 38.150 ;
        RECT 0.965 33.700 75.000 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 75.000 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 75.000 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 75.000 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 75.000 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 75.000 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 168.730 75.000 197.965 ;
        RECT 0.000 98.265 8.670 168.730 ;
        RECT 66.270 98.265 75.000 168.730 ;
        RECT 0.000 94.550 75.000 98.265 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vccd_lvc_clamped_pad

#--------EOF---------

MACRO sky130_ef_io__vccd_lvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vccd_lvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 -0.035 36.880 20.185 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 -0.035 49.255 22.865 ;
    END
  END DRN_LVC2
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 -0.035 20.495 1.450 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 -0.035 74.700 3.625 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 -0.035 44.440 0.290 ;
    END
  END BDY2_B2B
  PIN VCCD_PAD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 10.270 99.865 64.670 167.130 ;
    END
  END VCCD_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 6.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 6.865 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 74.785 197.805 ;
        RECT 16.655 -0.035 25.635 0.000 ;
        POLYGON 25.635 0.000 25.670 0.000 25.635 -0.035 ;
        RECT 26.210 -0.035 27.700 0.000 ;
        POLYGON 28.235 0.000 28.270 0.000 28.270 -0.035 ;
        RECT 28.270 -0.035 56.565 0.000 ;
      LAYER met2 ;
        RECT 0.490 3.905 74.700 194.395 ;
        RECT 0.490 3.625 54.435 3.905 ;
        RECT 0.490 1.730 54.715 3.625 ;
        RECT 20.775 0.570 54.715 1.730 ;
        RECT 20.775 0.005 34.160 0.570 ;
        RECT 44.720 0.005 54.715 0.570 ;
        RECT 20.775 0.000 34.440 0.005 ;
        RECT 20.925 -0.035 34.440 0.000 ;
        RECT 44.440 0.000 54.715 0.005 ;
        RECT 44.440 -0.035 53.535 0.000 ;
        RECT 54.095 -0.035 54.715 0.000 ;
      LAYER met3 ;
        RECT 0.490 23.265 74.700 189.480 ;
        RECT 0.490 20.585 37.980 23.265 ;
        RECT 0.490 7.265 25.600 20.585 ;
        RECT 24.900 0.000 25.600 7.265 ;
        RECT 37.280 0.000 37.980 20.585 ;
        RECT 49.655 7.265 74.700 23.265 ;
        RECT 49.655 0.000 50.355 7.265 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 168.730 75.000 197.965 ;
        RECT 0.000 98.265 8.670 168.730 ;
        RECT 66.270 98.265 75.000 168.730 ;
        RECT 0.000 94.550 75.000 98.265 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vccd_lvc_pad

#--------EOF---------

MACRO sky130_ef_io__vdda_hvc_clamped_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vdda_hvc_clamped_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN VDDA_PAD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 7.050 103.085 67.890 163.910 ;
    END
  END VDDA_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 12.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 12.925 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.630 189.565 0.640 189.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.360 189.565 74.370 189.575 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER pwell ;
        RECT 3.495 -1.100 11.285 21.755 ;
      LAYER nwell ;
        RECT 11.860 -1.350 70.965 0.170 ;
      LAYER li1 ;
        RECT 0.610 0.000 72.855 197.660 ;
        RECT 0.610 -0.970 11.155 0.000 ;
        RECT 12.035 -0.115 13.045 0.000 ;
        RECT 69.730 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met1 ;
        RECT 0.185 0.000 72.915 197.690 ;
        RECT 3.625 -0.905 8.855 0.000 ;
        RECT 12.035 -0.115 13.350 0.000 ;
        POLYGON 13.350 0.000 13.465 -0.115 13.350 -0.115 ;
        POLYGON 69.540 0.000 69.540 -0.115 69.425 -0.115 ;
        RECT 69.540 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met2 ;
        RECT 0.265 0.000 74.290 193.040 ;
        RECT 0.495 -2.035 24.395 0.000 ;
        RECT 25.895 -2.035 27.895 -0.115 ;
        RECT 50.390 -2.035 74.290 0.000 ;
      LAYER met3 ;
        RECT 0.240 13.325 74.290 197.965 ;
        RECT 24.795 0.000 49.990 13.325 ;
        RECT 25.895 -2.035 36.895 0.000 ;
        RECT 37.890 -2.035 48.890 0.000 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 165.510 75.000 197.965 ;
        RECT 0.000 101.485 5.450 165.510 ;
        RECT 69.490 101.485 75.000 165.510 ;
        RECT 0.000 94.550 75.000 101.485 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vdda_hvc_clamped_pad

#--------EOF---------

MACRO sky130_ef_io__vdda_hvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vdda_hvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.730 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.610 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 50.390 -2.035 74.290 23.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 -2.035 48.890 9.295 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.495 -2.035 24.395 0.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895 -2.035 36.895 0.690 ;
    END
  END SRC_BDY_HVC
  PIN VDDA_PAD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 7.050 103.085 67.890 163.910 ;
    END
  END VDDA_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.070 75.000 56.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 14.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 14.925 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 199.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 199.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.630 189.565 0.640 189.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.360 189.565 74.370 189.575 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER pwell ;
        RECT 3.495 -1.100 11.285 21.755 ;
      LAYER nwell ;
        RECT 11.860 -1.350 70.965 0.170 ;
      LAYER li1 ;
        RECT 0.610 0.000 72.855 197.660 ;
        RECT 0.610 -0.970 11.155 0.000 ;
        RECT 12.035 -0.115 13.045 0.000 ;
        RECT 69.730 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met1 ;
        RECT 0.185 0.000 72.915 197.690 ;
        RECT 3.625 -0.905 8.855 0.000 ;
        RECT 12.035 -0.115 13.350 0.000 ;
        POLYGON 13.350 0.000 13.465 -0.115 13.350 -0.115 ;
        POLYGON 69.540 0.000 69.540 -0.115 69.425 -0.115 ;
        RECT 69.540 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met2 ;
        RECT 0.265 23.905 74.290 193.040 ;
        RECT 0.265 0.300 50.110 23.905 ;
        RECT 24.675 0.000 50.110 0.300 ;
        RECT 25.895 -2.035 27.895 -0.115 ;
      LAYER met3 ;
        RECT 0.240 15.325 74.290 197.965 ;
        RECT 24.795 9.695 49.990 15.325 ;
        RECT 24.795 1.090 37.490 9.695 ;
        RECT 24.795 0.690 25.495 1.090 ;
        RECT 37.295 0.690 37.490 1.090 ;
        RECT 49.290 0.690 49.990 9.695 ;
      LAYER met4 ;
        RECT 1.205 197.965 74.225 199.965 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.000 93.145 75.000 173.350 ;
        RECT 0.000 92.965 0.715 93.145 ;
        RECT 0.000 67.600 0.715 68.000 ;
        RECT 1.670 67.600 73.330 93.145 ;
        RECT 0.000 66.500 75.000 67.600 ;
        RECT 0.000 61.650 0.715 62.050 ;
        RECT 1.670 61.650 73.330 66.500 ;
        RECT 0.000 60.650 75.000 61.650 ;
        RECT 1.670 56.470 73.330 60.650 ;
        RECT 1.670 51.090 73.330 53.670 ;
        RECT 0.000 50.790 75.000 51.090 ;
        RECT 1.670 50.010 73.330 50.790 ;
        RECT 0.000 46.030 75.000 46.200 ;
        RECT 0.000 45.300 0.715 45.700 ;
        RECT 1.670 45.300 73.330 45.930 ;
        RECT 0.000 44.200 75.000 45.300 ;
        RECT 0.000 39.150 0.715 39.550 ;
        RECT 1.670 39.150 73.330 44.200 ;
        RECT 0.000 38.150 75.000 39.150 ;
        RECT 0.000 34.300 0.715 34.700 ;
        RECT 1.670 34.300 73.330 38.150 ;
        RECT 0.000 33.300 75.000 34.300 ;
        RECT 0.000 29.450 0.715 29.850 ;
        RECT 1.670 29.450 73.330 33.300 ;
        RECT 0.000 28.450 75.000 29.450 ;
        RECT 0.000 23.400 0.715 23.800 ;
        RECT 1.670 23.400 73.330 28.450 ;
        RECT 0.000 22.400 75.000 23.400 ;
        RECT 0.000 17.565 0.525 17.750 ;
        RECT 0.000 17.445 0.715 17.565 ;
        RECT 0.000 17.350 0.525 17.445 ;
        RECT 1.670 17.350 73.330 22.400 ;
        RECT 0.000 16.750 75.000 17.350 ;
        RECT 0.000 16.685 0.525 16.750 ;
        RECT 1.365 16.685 73.635 16.750 ;
        RECT 0.000 16.565 75.000 16.685 ;
        RECT 0.000 16.350 0.525 16.565 ;
        RECT 0.000 12.500 0.715 12.900 ;
        RECT 1.365 12.500 73.635 16.565 ;
        RECT 0.000 11.500 75.000 12.500 ;
        RECT 0.000 6.450 0.715 6.850 ;
        RECT 1.670 6.450 73.330 11.500 ;
        RECT 0.000 5.450 75.000 6.450 ;
        RECT 1.670 0.000 73.330 5.450 ;
      LAYER met5 ;
        RECT 0.000 165.510 75.000 199.965 ;
        RECT 0.000 101.485 5.450 165.510 ;
        RECT 69.490 101.485 75.000 165.510 ;
        RECT 0.000 94.550 75.000 101.485 ;
        RECT 0.000 93.645 0.715 94.550 ;
        RECT 2.870 93.645 72.130 94.550 ;
        RECT 0.000 93.145 75.000 93.645 ;
        RECT 0.000 92.950 0.715 93.145 ;
        RECT 0.000 67.100 0.715 68.000 ;
        RECT 2.870 67.100 72.130 93.145 ;
        RECT 0.000 66.400 75.000 67.100 ;
        RECT 0.000 61.250 0.715 62.150 ;
        RECT 2.870 61.250 72.130 66.400 ;
        RECT 0.000 60.550 75.000 61.250 ;
        RECT 2.870 56.300 72.130 60.550 ;
        RECT 0.000 54.700 75.000 56.300 ;
        RECT 0.000 44.800 0.715 45.700 ;
        RECT 2.870 44.800 72.130 54.700 ;
        RECT 0.000 44.100 75.000 44.800 ;
        RECT 0.000 38.750 0.715 39.650 ;
        RECT 2.870 38.750 72.130 44.100 ;
        RECT 0.000 38.100 75.000 38.750 ;
        RECT 0.000 38.050 0.715 38.100 ;
        RECT 0.000 33.900 0.715 34.805 ;
        RECT 2.870 33.900 72.130 38.100 ;
        RECT 0.000 33.250 75.000 33.900 ;
        RECT 0.000 33.200 0.715 33.250 ;
        RECT 0.000 29.050 0.715 29.950 ;
        RECT 2.870 29.050 72.130 33.250 ;
        RECT 0.000 28.350 75.000 29.050 ;
        RECT 0.000 23.000 0.715 23.900 ;
        RECT 2.870 23.000 72.130 28.350 ;
        RECT 0.000 22.300 75.000 23.000 ;
        RECT 0.000 16.950 0.715 17.850 ;
        RECT 2.870 16.950 72.130 22.300 ;
        RECT 0.000 16.300 75.000 16.950 ;
        RECT 0.000 16.250 0.715 16.300 ;
        RECT 2.870 16.250 72.130 16.300 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 0.000 12.100 0.715 13.000 ;
        RECT 2.870 12.100 72.130 13.000 ;
        RECT 0.000 11.400 75.000 12.100 ;
        RECT 0.000 6.045 0.715 6.950 ;
        RECT 2.870 6.045 72.130 11.400 ;
        RECT 0.000 5.350 75.000 6.045 ;
        RECT 2.870 0.100 72.130 5.350 ;
  END
END sky130_ef_io__vdda_hvc_pad

#--------EOF---------

MACRO sky130_ef_io__vdda_lvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vdda_lvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 -0.035 36.880 20.185 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 -0.035 49.255 22.865 ;
    END
  END DRN_LVC2
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 -0.035 20.495 1.450 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 -0.035 74.700 3.625 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 -0.035 44.440 0.290 ;
    END
  END BDY2_B2B
  PIN VDDA_PAD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 10.270 99.865 64.670 167.130 ;
    END
  END VDDA_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 12.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 12.925 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 74.785 197.805 ;
        RECT 16.655 -0.035 25.635 0.000 ;
        POLYGON 25.635 0.000 25.670 0.000 25.635 -0.035 ;
        RECT 26.210 -0.035 27.700 0.000 ;
        POLYGON 28.235 0.000 28.270 0.000 28.270 -0.035 ;
        RECT 28.270 -0.035 56.565 0.000 ;
      LAYER met2 ;
        RECT 0.490 3.905 74.700 194.395 ;
        RECT 0.490 3.625 54.435 3.905 ;
        RECT 0.490 1.730 54.715 3.625 ;
        RECT 20.775 0.570 54.715 1.730 ;
        RECT 20.775 0.005 34.160 0.570 ;
        RECT 44.720 0.005 54.715 0.570 ;
        RECT 20.775 0.000 34.440 0.005 ;
        RECT 20.925 -0.035 34.440 0.000 ;
        RECT 44.440 0.000 54.715 0.005 ;
        RECT 44.440 -0.035 53.535 0.000 ;
        RECT 54.095 -0.035 54.715 0.000 ;
      LAYER met3 ;
        RECT 0.490 23.265 74.700 189.480 ;
        RECT 0.490 20.585 37.980 23.265 ;
        RECT 0.490 13.325 25.600 20.585 ;
        RECT 24.900 0.000 25.600 13.325 ;
        RECT 37.280 0.000 37.980 20.585 ;
        RECT 49.655 13.325 74.700 23.265 ;
        RECT 49.655 0.000 50.355 13.325 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 168.730 75.000 197.965 ;
        RECT 0.000 98.265 8.670 168.730 ;
        RECT 66.270 98.265 75.000 168.730 ;
        RECT 0.000 94.550 75.000 98.265 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vdda_lvc_pad

#--------EOF---------

MACRO sky130_ef_io__vddio_hvc_clamped_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vddio_hvc_clamped_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN VDDIO_PAD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 7.050 103.085 67.890 163.910 ;
    END
  END VDDIO_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 17.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 17.765 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER pwell ;
        RECT 3.495 -1.100 11.285 21.755 ;
      LAYER nwell ;
        RECT 11.860 -1.350 70.965 0.170 ;
      LAYER li1 ;
        RECT 0.610 0.000 72.855 197.660 ;
        RECT 0.610 -0.970 11.155 0.000 ;
        RECT 12.035 -0.115 13.045 0.000 ;
        RECT 69.730 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met1 ;
        RECT 0.185 0.000 72.915 197.690 ;
        RECT 3.625 -0.905 8.855 0.000 ;
        RECT 12.035 -0.115 13.350 0.000 ;
        POLYGON 13.350 0.000 13.465 -0.115 13.350 -0.115 ;
        POLYGON 69.540 0.000 69.540 -0.115 69.425 -0.115 ;
        RECT 69.540 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met2 ;
        RECT 0.265 0.000 74.290 193.040 ;
        RECT 0.495 -2.035 24.395 0.000 ;
        RECT 25.895 -2.035 27.895 -0.115 ;
        RECT 50.390 -2.035 74.290 0.000 ;
      LAYER met3 ;
        RECT 0.240 18.165 74.290 197.965 ;
        RECT 24.795 0.000 49.990 18.165 ;
        RECT 25.895 -2.035 36.895 0.000 ;
        RECT 37.890 -2.035 48.890 0.000 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 165.510 75.000 197.965 ;
        RECT 0.000 101.485 5.450 165.510 ;
        RECT 69.490 101.485 75.000 165.510 ;
        RECT 0.000 94.550 75.000 101.485 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vddio_hvc_clamped_pad

#--------EOF---------

MACRO sky130_ef_io__vddio_hvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vddio_hvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 50.390 -2.035 74.290 23.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 -2.035 48.890 9.295 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.495 -2.035 24.395 0.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895 -2.035 36.895 0.690 ;
    END
  END SRC_BDY_HVC
  PIN VDDIO_PAD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 7.050 103.085 67.890 163.910 ;
    END
  END VDDIO_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 17.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 17.765 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER pwell ;
        RECT 3.495 -1.100 11.285 21.755 ;
      LAYER nwell ;
        RECT 11.860 -1.350 70.965 0.170 ;
      LAYER li1 ;
        RECT 0.610 0.000 72.855 197.660 ;
        RECT 0.610 -0.970 11.155 0.000 ;
        RECT 12.035 -0.115 13.045 0.000 ;
        RECT 69.730 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met1 ;
        RECT 0.185 0.000 72.915 197.690 ;
        RECT 3.625 -0.905 8.855 0.000 ;
        RECT 12.035 -0.115 13.350 0.000 ;
        POLYGON 13.350 0.000 13.465 -0.115 13.350 -0.115 ;
        POLYGON 69.540 0.000 69.540 -0.115 69.425 -0.115 ;
        RECT 69.540 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met2 ;
        RECT 0.265 23.905 74.290 193.040 ;
        RECT 0.265 0.300 50.110 23.905 ;
        RECT 24.675 0.000 50.110 0.300 ;
        RECT 25.895 -2.035 27.895 -0.115 ;
      LAYER met3 ;
        RECT 0.240 18.165 74.290 197.965 ;
        RECT 24.795 9.695 49.990 18.165 ;
        RECT 24.795 1.090 37.490 9.695 ;
        RECT 24.795 0.690 25.495 1.090 ;
        RECT 37.295 0.690 37.490 1.090 ;
        RECT 49.290 0.690 49.990 9.695 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 165.510 75.000 197.965 ;
        RECT 0.000 101.485 5.450 165.510 ;
        RECT 69.490 101.485 75.000 165.510 ;
        RECT 0.000 94.550 75.000 101.485 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vddio_hvc_pad

#--------EOF---------

MACRO sky130_ef_io__vddio_lvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vddio_lvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 -0.035 36.880 20.185 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 -0.035 49.255 22.865 ;
    END
  END DRN_LVC2
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 -0.035 20.495 1.450 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 -0.035 74.700 3.625 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 -0.035 44.440 0.290 ;
    END
  END BDY2_B2B
  PIN VDDIO_PAD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 10.270 99.865 64.670 167.130 ;
    END
  END VDDIO_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 17.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 17.765 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 74.785 197.805 ;
        RECT 16.655 -0.035 25.635 0.000 ;
        POLYGON 25.635 0.000 25.670 0.000 25.635 -0.035 ;
        RECT 26.210 -0.035 27.700 0.000 ;
        POLYGON 28.235 0.000 28.270 0.000 28.270 -0.035 ;
        RECT 28.270 -0.035 56.565 0.000 ;
      LAYER met2 ;
        RECT 0.490 3.905 74.700 194.395 ;
        RECT 0.490 3.625 54.435 3.905 ;
        RECT 0.490 1.730 54.715 3.625 ;
        RECT 20.775 0.570 54.715 1.730 ;
        RECT 20.775 0.005 34.160 0.570 ;
        RECT 44.720 0.005 54.715 0.570 ;
        RECT 20.775 0.000 34.440 0.005 ;
        RECT 20.925 -0.035 34.440 0.000 ;
        RECT 44.440 0.000 54.715 0.005 ;
        RECT 44.440 -0.035 53.535 0.000 ;
        RECT 54.095 -0.035 54.715 0.000 ;
      LAYER met3 ;
        RECT 0.490 23.265 74.700 189.480 ;
        RECT 0.490 20.585 37.980 23.265 ;
        RECT 0.490 18.165 25.600 20.585 ;
        RECT 24.900 0.000 25.600 18.165 ;
        RECT 37.280 0.000 37.980 20.585 ;
        RECT 49.655 18.165 74.700 23.265 ;
        RECT 49.655 0.000 50.355 18.165 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 168.730 75.000 197.965 ;
        RECT 0.000 98.265 8.670 168.730 ;
        RECT 66.270 98.265 75.000 168.730 ;
        RECT 0.000 94.550 75.000 98.265 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vddio_lvc_pad

#--------EOF---------

MACRO sky130_ef_io__vssa_hvc_clamped_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssa_hvc_clamped_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSA_PAD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 7.050 103.085 67.890 163.910 ;
    END
  END VSSA_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 30.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 34.725 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.360 189.565 74.370 189.575 ;
    END
  END VSSIO
  OBS
      LAYER nwell ;
        RECT 11.860 -1.350 70.965 0.170 ;
      LAYER li1 ;
        RECT 1.070 0.000 72.775 197.660 ;
        RECT 12.065 -0.145 13.045 0.000 ;
        RECT 69.760 -0.145 70.650 0.000 ;
        RECT 12.065 -1.035 70.650 -0.145 ;
      LAYER met1 ;
        RECT 0.185 0.000 73.620 197.690 ;
        RECT 12.035 -0.115 13.350 0.000 ;
        POLYGON 13.350 0.000 13.465 -0.115 13.350 -0.115 ;
        POLYGON 69.540 0.000 69.540 -0.115 69.425 -0.115 ;
        RECT 69.540 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met2 ;
        RECT 0.265 0.000 74.290 193.040 ;
        RECT 0.495 -2.035 24.395 0.000 ;
        RECT 25.895 -2.035 27.895 -0.115 ;
        RECT 50.390 -2.035 74.290 0.000 ;
      LAYER met3 ;
        RECT 0.240 35.125 74.290 193.065 ;
        RECT 0.240 30.880 49.990 35.125 ;
        RECT 24.795 0.000 49.990 30.880 ;
        RECT 25.895 -2.035 36.895 0.000 ;
        RECT 37.890 -2.035 48.890 0.000 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 54.470 73.330 55.100 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 1.670 45.300 73.330 45.930 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 165.510 75.000 197.965 ;
        RECT 0.000 101.485 5.450 165.510 ;
        RECT 69.490 101.485 75.000 165.510 ;
        RECT 0.000 94.550 75.000 101.485 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssa_hvc_clamped_pad

#--------EOF---------

MACRO sky130_ef_io__vssa_hvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssa_hvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 50.390 -2.035 74.290 23.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 -2.035 48.890 10.345 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.495 -2.035 24.395 0.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895 -2.035 36.895 10.390 ;
    END
  END SRC_BDY_HVC
  PIN VSSA_PAD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 7.050 103.085 67.890 163.910 ;
    END
  END VSSA_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 30.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 34.725 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.360 189.565 74.370 189.575 ;
    END
  END VSSIO
  OBS
      LAYER nwell ;
        RECT 11.860 -1.350 70.965 0.170 ;
      LAYER li1 ;
        RECT 1.070 0.000 72.775 197.660 ;
        RECT 12.065 -0.145 13.045 0.000 ;
        RECT 69.760 -0.145 70.650 0.000 ;
        RECT 12.065 -1.035 70.650 -0.145 ;
      LAYER met1 ;
        RECT 0.185 0.000 73.620 197.690 ;
        RECT 12.035 -0.115 13.350 0.000 ;
        POLYGON 13.350 0.000 13.465 -0.115 13.350 -0.115 ;
        POLYGON 69.540 0.000 69.540 -0.115 69.425 -0.115 ;
        RECT 69.540 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met2 ;
        RECT 0.265 23.905 74.290 193.040 ;
        RECT 0.265 0.300 50.110 23.905 ;
        RECT 24.675 0.000 50.110 0.300 ;
        RECT 25.895 -2.035 27.895 -0.115 ;
      LAYER met3 ;
        RECT 0.240 35.125 74.290 193.065 ;
        RECT 0.240 30.880 49.990 35.125 ;
        RECT 24.795 10.790 49.990 30.880 ;
        RECT 24.795 10.345 25.495 10.790 ;
        RECT 37.295 10.745 49.990 10.790 ;
        RECT 37.295 10.345 37.490 10.745 ;
        RECT 49.290 10.345 49.990 10.745 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 54.470 73.330 55.100 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 1.670 45.300 73.330 45.930 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 165.510 75.000 197.965 ;
        RECT 0.000 101.485 5.450 165.510 ;
        RECT 69.490 101.485 75.000 165.510 ;
        RECT 0.000 94.550 75.000 101.485 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssa_hvc_pad

#--------EOF---------

MACRO sky130_ef_io__vssa_lvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssa_lvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.090 75.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 46.330 75.000 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 -0.035 36.880 20.185 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 -0.035 49.255 22.865 ;
    END
  END DRN_LVC2
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 -0.035 20.495 1.450 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 -0.035 74.700 3.625 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 -0.035 44.440 0.290 ;
    END
  END BDY2_B2B
  PIN VSSA_PAD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 10.270 99.865 64.670 167.130 ;
    END
  END VSSA_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 34.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 34.725 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 74.785 197.805 ;
        RECT 16.655 -0.035 25.635 0.000 ;
        POLYGON 25.635 0.000 25.670 0.000 25.635 -0.035 ;
        RECT 26.210 -0.035 27.700 0.000 ;
        POLYGON 28.235 0.000 28.270 0.000 28.270 -0.035 ;
        RECT 28.270 -0.035 56.565 0.000 ;
      LAYER met2 ;
        RECT 0.500 3.905 74.700 194.395 ;
        RECT 0.500 3.625 54.435 3.905 ;
        RECT 0.500 1.730 54.715 3.625 ;
        RECT 20.775 0.570 54.715 1.730 ;
        RECT 20.775 0.005 34.160 0.570 ;
        RECT 44.720 0.005 54.715 0.570 ;
        RECT 20.775 0.000 34.440 0.005 ;
        RECT 20.925 -0.035 34.440 0.000 ;
        RECT 44.440 0.000 54.715 0.005 ;
        RECT 44.440 -0.035 53.535 0.000 ;
        RECT 54.095 -0.035 54.715 0.000 ;
      LAYER met3 ;
        RECT 0.490 35.125 74.700 189.480 ;
        RECT 24.900 23.265 50.355 35.125 ;
        RECT 24.900 20.585 37.980 23.265 ;
        RECT 24.900 1.545 25.600 20.585 ;
        RECT 37.280 1.545 37.980 20.585 ;
        RECT 49.655 1.545 50.355 23.265 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 168.730 75.000 197.965 ;
        RECT 0.000 98.265 8.670 168.730 ;
        RECT 66.270 98.265 75.000 168.730 ;
        RECT 0.000 94.550 75.000 98.265 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssa_lvc_pad

#--------EOF---------

MACRO sky130_ef_io__vssd_hvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssd_hvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 50.390 -2.035 74.290 23.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 -2.035 48.890 10.345 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.495 -2.035 24.395 0.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895 -2.035 36.895 10.390 ;
    END
  END SRC_BDY_HVC
  PIN VSSD_PAD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 7.050 103.085 67.890 163.910 ;
    END
  END VSSD_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 30.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 39.565 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER nwell ;
        RECT 11.860 -1.350 70.965 0.170 ;
      LAYER li1 ;
        RECT 1.070 0.000 72.775 197.660 ;
        RECT 12.065 -0.145 13.045 0.000 ;
        RECT 69.760 -0.145 70.650 0.000 ;
        RECT 12.065 -1.035 70.650 -0.145 ;
      LAYER met1 ;
        RECT 0.185 0.000 73.620 197.690 ;
        RECT 12.035 -0.115 13.350 0.000 ;
        POLYGON 13.350 0.000 13.465 -0.115 13.350 -0.115 ;
        POLYGON 69.540 0.000 69.540 -0.115 69.425 -0.115 ;
        RECT 69.540 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met2 ;
        RECT 0.265 23.905 74.290 193.040 ;
        RECT 0.265 0.300 50.110 23.905 ;
        RECT 24.675 0.000 50.110 0.300 ;
        RECT 25.895 -2.035 27.895 -0.115 ;
      LAYER met3 ;
        RECT 0.240 39.965 74.290 193.065 ;
        RECT 0.240 30.880 49.990 39.965 ;
        RECT 24.795 10.790 49.990 30.880 ;
        RECT 24.795 10.345 25.495 10.790 ;
        RECT 37.295 10.745 49.990 10.790 ;
        RECT 37.295 10.345 37.490 10.745 ;
        RECT 49.290 10.345 49.990 10.745 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 165.510 75.000 197.965 ;
        RECT 0.000 101.485 5.450 165.510 ;
        RECT 69.490 101.485 75.000 165.510 ;
        RECT 0.000 94.550 75.000 101.485 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssd_hvc_pad

#--------EOF---------

MACRO sky130_ef_io__vssd_lvc_clamped2_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssd_lvc_clamped2_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSD_PAD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 10.270 99.865 64.670 167.130 ;
    END
  END VSSD_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 76.470 197.930 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 39.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 39.565 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 75.000 197.805 ;
        RECT 16.655 -0.035 56.565 0.000 ;
        RECT 20.925 -0.815 56.565 -0.035 ;
        RECT 76.200 -0.815 85.935 75.350 ;
        RECT 20.925 -6.920 85.935 -0.815 ;
        RECT 20.925 -10.920 81.935 -6.920 ;
        POLYGON 81.935 -6.920 85.935 -6.920 81.935 -10.920 ;
      LAYER met2 ;
        RECT 0.000 44.200 75.000 197.930 ;
        RECT 76.200 46.560 85.935 197.930 ;
        RECT 0.000 44.165 86.140 44.200 ;
        RECT -10.975 39.550 86.140 44.165 ;
        RECT -10.975 39.515 75.000 39.550 ;
        RECT 0.000 0.000 75.000 39.515 ;
        RECT 76.200 23.390 85.935 37.800 ;
        RECT 0.500 -0.035 20.495 0.000 ;
        RECT 20.925 -0.035 53.535 0.000 ;
        RECT 54.095 -0.035 74.700 0.000 ;
      LAYER met3 ;
        RECT -10.975 39.515 -0.895 44.165 ;
        RECT 0.000 39.965 75.000 197.930 ;
        RECT 76.200 173.715 85.935 197.930 ;
        RECT 0.000 0.000 0.100 39.965 ;
        RECT 24.900 0.000 50.355 39.965 ;
        RECT 75.605 39.550 86.140 44.200 ;
        RECT 76.200 23.765 85.935 28.415 ;
        RECT 26.000 -0.035 36.880 0.000 ;
        RECT 38.380 -0.035 49.255 0.000 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 76.470 173.750 85.935 197.930 ;
        RECT 74.785 173.715 85.935 173.750 ;
        RECT 0.000 93.365 75.000 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.000 66.900 75.000 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.000 61.050 75.000 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.000 55.100 75.000 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.000 44.600 75.000 45.300 ;
        RECT -10.975 39.550 0.000 44.165 ;
        RECT -10.975 39.515 0.070 39.550 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 75.000 39.550 86.140 44.200 ;
        RECT 0.000 38.550 75.000 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.000 33.700 75.000 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.000 28.850 75.000 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 75.000 23.800 85.935 28.415 ;
        RECT 74.935 23.765 85.935 23.800 ;
        RECT 0.000 22.800 75.000 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.000 16.750 75.000 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.000 11.900 75.000 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.000 5.850 75.000 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 168.730 75.000 197.965 ;
        RECT 0.000 98.265 8.670 168.730 ;
        RECT 66.270 98.265 75.000 168.730 ;
        RECT 0.000 94.550 75.000 98.265 ;
        RECT 2.870 16.250 72.130 94.550 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssd_lvc_clamped2_pad

#--------EOF---------

MACRO sky130_ef_io__vssd_lvc_clamped3_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssd_lvc_clamped3_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSD_PAD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 10.270 99.865 64.670 167.130 ;
    END
  END VSSD_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 76.470 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  PIN VSSD1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER met3 ;
        RECT 0.500 -9.480 24.500 26.400 ;
    END
    PORT
      CLASS CORE ;
      LAYER met3 ;
        RECT 50.755 -9.510 74.700 27.120 ;
    END
  END VSSD1
  PIN VCCD1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER met3 ;
        RECT 26.000 -9.490 49.255 -2.290 ;
    END
  END VCCD1
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 75.000 197.805 ;
        RECT 16.655 -0.035 56.565 0.000 ;
        RECT 20.925 -0.780 56.565 -0.035 ;
        RECT 76.200 -0.780 85.935 75.385 ;
        RECT 20.925 -6.885 85.935 -0.780 ;
        RECT 20.925 -10.885 81.935 -6.885 ;
        POLYGON 81.935 -6.885 85.935 -6.885 81.935 -10.885 ;
      LAYER met2 ;
        RECT 0.500 0.000 75.000 197.965 ;
        RECT 76.200 23.425 85.935 197.965 ;
        RECT 0.500 -0.035 20.495 0.000 ;
        RECT 20.925 -0.035 53.535 0.000 ;
        RECT 54.095 -0.035 74.700 0.000 ;
      LAYER met3 ;
        RECT 0.500 27.520 75.000 197.965 ;
        RECT 76.200 173.750 85.935 197.965 ;
        RECT 0.500 26.800 50.355 27.520 ;
        RECT 24.900 0.000 50.355 26.800 ;
        RECT 76.200 23.800 85.935 28.450 ;
        RECT 26.000 -2.290 36.880 0.000 ;
        RECT 38.380 -2.290 49.255 0.000 ;
      LAYER met4 ;
        RECT 1.605 173.350 73.825 197.965 ;
        RECT 76.470 173.750 85.935 197.965 ;
        RECT 0.965 93.365 75.000 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 75.000 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 75.000 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 75.000 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 75.000 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 75.000 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 75.000 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 75.000 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 75.000 23.800 85.935 28.450 ;
        RECT 0.965 22.800 75.000 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 75.000 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 75.000 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 75.000 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 168.730 75.000 197.965 ;
        RECT 0.000 98.265 8.670 168.730 ;
        RECT 66.270 98.265 75.000 168.730 ;
        RECT 0.000 94.550 75.000 98.265 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssd_lvc_clamped3_pad

#--------EOF---------

MACRO sky130_ef_io__vssd_lvc_clamped_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssd_lvc_clamped_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSD_PAD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 10.270 99.865 64.670 167.130 ;
    END
  END VSSD_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 0.705 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 39.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 39.565 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 75.000 197.805 ;
        RECT 75.245 34.455 86.195 38.325 ;
        RECT 16.655 -0.035 56.565 0.000 ;
        RECT 20.495 -0.815 56.565 -0.035 ;
        RECT 76.200 -0.815 85.935 34.455 ;
        RECT 20.495 -1.015 85.935 -0.815 ;
        POLYGON 18.655 -1.015 18.655 -3.015 16.655 -3.015 ;
        RECT 18.655 -3.015 85.935 -1.015 ;
        RECT 16.655 -6.535 85.935 -3.015 ;
        RECT 16.655 -8.535 81.935 -6.535 ;
        POLYGON 16.655 -8.535 18.655 -8.535 18.655 -10.535 ;
        RECT 18.655 -10.535 81.935 -8.535 ;
        POLYGON 81.935 -6.535 85.935 -6.535 81.935 -10.535 ;
      LAYER met2 ;
        RECT 0.500 44.200 75.000 194.395 ;
        RECT 0.500 39.550 86.140 44.200 ;
        RECT 0.500 0.000 75.000 39.550 ;
        RECT 75.245 34.455 86.195 38.325 ;
        RECT 0.500 -0.035 20.495 0.000 ;
        RECT 20.925 -0.035 53.535 0.000 ;
        RECT 54.095 -0.035 74.700 0.000 ;
      LAYER met3 ;
        RECT 0.500 39.965 75.000 193.570 ;
        RECT 24.900 0.000 50.355 39.965 ;
        RECT 75.605 39.550 86.140 44.200 ;
        RECT 75.440 34.695 86.140 38.160 ;
        RECT 26.000 -0.035 36.880 0.000 ;
        RECT 38.380 -0.035 49.255 0.000 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 75.000 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 75.000 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 75.000 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 75.000 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 75.000 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 75.000 39.550 86.140 44.200 ;
        RECT 0.965 38.550 75.000 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 75.000 34.700 86.165 38.150 ;
        RECT 0.965 33.700 75.000 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 75.000 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 75.000 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 75.000 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 75.000 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 75.000 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 168.730 75.000 197.965 ;
        RECT 0.000 98.265 8.670 168.730 ;
        RECT 66.270 98.265 75.000 168.730 ;
        RECT 0.000 94.550 75.000 98.265 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssd_lvc_clamped_pad

#--------EOF---------

MACRO sky130_ef_io__vssd_lvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssd_lvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 -0.035 36.880 20.185 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 -0.035 49.255 22.865 ;
    END
  END DRN_LVC2
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 -0.035 20.495 1.450 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 -0.035 74.700 3.625 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 -0.035 44.440 0.290 ;
    END
  END BDY2_B2B
  PIN VSSD_PAD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 10.270 99.865 64.670 167.130 ;
    END
  END VSSD_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.225 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.205 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 39.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 39.565 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 74.785 197.805 ;
        RECT 16.655 -0.035 25.635 0.000 ;
        POLYGON 25.635 0.000 25.670 0.000 25.635 -0.035 ;
        RECT 26.210 -0.035 27.700 0.000 ;
        POLYGON 28.235 0.000 28.270 0.000 28.270 -0.035 ;
        RECT 28.270 -0.035 56.565 0.000 ;
      LAYER met2 ;
        RECT 0.500 3.905 74.700 194.395 ;
        RECT 0.500 3.625 54.435 3.905 ;
        RECT 0.500 1.730 54.715 3.625 ;
        RECT 20.775 0.570 54.715 1.730 ;
        RECT 20.775 0.005 34.160 0.570 ;
        RECT 44.720 0.005 54.715 0.570 ;
        RECT 20.775 0.000 34.440 0.005 ;
        RECT 20.925 -0.035 34.440 0.000 ;
        RECT 44.440 0.000 54.715 0.005 ;
        RECT 44.440 -0.035 53.535 0.000 ;
        RECT 54.095 -0.035 54.715 0.000 ;
      LAYER met3 ;
        RECT 0.500 39.965 74.700 189.480 ;
        RECT 24.900 23.265 50.355 39.965 ;
        RECT 24.900 20.585 37.980 23.265 ;
        RECT 24.900 17.755 25.600 20.585 ;
        RECT 37.280 17.755 37.980 20.585 ;
        RECT 49.655 17.755 50.355 23.265 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 168.730 75.000 197.965 ;
        RECT 0.000 98.265 8.670 168.730 ;
        RECT 66.270 98.265 75.000 168.730 ;
        RECT 0.000 94.550 75.000 98.265 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssd_lvc_pad

#--------EOF---------

MACRO sky130_ef_io__vssio_hvc_clamped_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssio_hvc_clamped_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSIO_PAD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 7.050 103.085 67.890 163.910 ;
    END
  END VSSIO_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.630 189.565 0.640 189.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.250 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 23.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 23.815 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER nwell ;
        RECT 11.860 -1.350 70.965 0.170 ;
      LAYER li1 ;
        RECT 1.070 0.000 72.775 197.660 ;
        RECT 12.065 -0.145 13.045 0.000 ;
        RECT 69.760 -0.145 70.650 0.000 ;
        RECT 12.065 -1.035 70.650 -0.145 ;
      LAYER met1 ;
        RECT 0.185 0.000 73.620 197.690 ;
        RECT 12.035 -0.115 13.350 0.000 ;
        POLYGON 13.350 0.000 13.465 -0.115 13.350 -0.115 ;
        POLYGON 69.540 0.000 69.540 -0.115 69.425 -0.115 ;
        RECT 69.540 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met2 ;
        RECT 0.265 0.000 74.290 193.040 ;
        RECT 0.495 -2.035 24.395 0.000 ;
        RECT 25.895 -2.035 27.895 -0.115 ;
        RECT 50.390 -2.035 74.290 0.000 ;
      LAYER met3 ;
        RECT 0.240 24.215 74.290 197.965 ;
        RECT 24.795 0.000 49.990 24.215 ;
        RECT 25.895 -2.035 36.895 0.000 ;
        RECT 37.890 -2.035 48.890 0.000 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 165.510 75.000 197.965 ;
        RECT 0.000 101.485 5.450 165.510 ;
        RECT 69.490 101.485 75.000 165.510 ;
        RECT 0.000 94.550 75.000 101.485 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssio_hvc_clamped_pad

#--------EOF---------

MACRO sky130_ef_io__vssio_hvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssio_hvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 50.390 -2.035 74.290 23.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 -2.035 48.890 10.345 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.495 -2.035 24.395 0.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895 -2.035 36.895 10.390 ;
    END
  END SRC_BDY_HVC
  PIN VSSIO_PAD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 7.050 103.085 67.890 163.910 ;
    END
  END VSSIO_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.630 189.565 0.640 189.575 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.250 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 -2.035 24.395 23.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 -2.035 74.290 23.815 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER nwell ;
        RECT 11.860 -1.350 70.965 0.170 ;
      LAYER li1 ;
        RECT 1.070 0.000 72.775 197.660 ;
        RECT 12.065 -0.145 13.045 0.000 ;
        RECT 69.760 -0.145 70.650 0.000 ;
        RECT 12.065 -1.035 70.650 -0.145 ;
      LAYER met1 ;
        RECT 0.185 0.000 73.620 197.690 ;
        RECT 12.035 -0.115 13.350 0.000 ;
        POLYGON 13.350 0.000 13.465 -0.115 13.350 -0.115 ;
        POLYGON 69.540 0.000 69.540 -0.115 69.425 -0.115 ;
        RECT 69.540 -0.115 70.680 0.000 ;
        RECT 12.035 -1.065 70.680 -0.115 ;
      LAYER met2 ;
        RECT 0.265 23.905 74.290 193.040 ;
        RECT 0.265 0.300 50.110 23.905 ;
        RECT 24.675 0.000 50.110 0.300 ;
        RECT 25.895 -2.035 27.895 -0.115 ;
      LAYER met3 ;
        RECT 0.240 24.215 74.290 197.965 ;
        RECT 24.795 10.790 49.990 24.215 ;
        RECT 24.795 10.345 25.495 10.790 ;
        RECT 37.295 10.745 49.990 10.790 ;
        RECT 37.295 10.345 37.490 10.745 ;
        RECT 49.290 10.345 49.990 10.745 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 165.510 75.000 197.965 ;
        RECT 0.000 101.485 5.450 165.510 ;
        RECT 69.490 101.485 75.000 165.510 ;
        RECT 0.000 94.550 75.000 101.485 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssio_hvc_pad

#--------EOF---------

MACRO sky130_ef_io__vssio_lvc_pad
  CLASS PAD POWER ;
  FOREIGN sky130_ef_io__vssio_lvc_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 75.000 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 1.270 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 75.000 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 1.270 49.310 ;
    END
  END AMUXBUS_B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 -0.035 36.880 20.185 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 -0.035 49.255 22.865 ;
    END
  END DRN_LVC2
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 -0.035 20.495 1.450 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 -0.035 74.700 3.625 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 -0.035 44.440 0.290 ;
    END
  END BDY2_B2B
  PIN VSSIO_PAD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 10.270 99.865 64.670 167.130 ;
    END
  END VSSIO_PAD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.700 75.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.805 75.000 38.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.610 75.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 75.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 75.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.700 75.000 38.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 1.270 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 1.270 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.000 75.000 16.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.900 75.000 16.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.950 75.000 33.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.850 75.000 33.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.150 75.000 66.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.050 75.000 66.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.100 75.000 5.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.000 75.000 5.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.000 75.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.850 75.000 22.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.750 75.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.000 75.000 92.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.950 75.000 11.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.850 75.000 11.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 50.755 -0.035 74.700 23.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 -0.035 24.500 23.815 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.900 75.000 28.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.800 75.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.750 75.000 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.650 75.000 44.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.550 75.000 44.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.300 75.000 60.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.200 75.000 60.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER li1 ;
        RECT 0.240 0.985 74.755 197.745 ;
      LAYER met1 ;
        RECT 0.120 0.000 74.785 197.805 ;
        RECT 16.655 -0.035 25.635 0.000 ;
        POLYGON 25.635 0.000 25.670 0.000 25.635 -0.035 ;
        RECT 26.210 -0.035 27.700 0.000 ;
        POLYGON 28.235 0.000 28.270 0.000 28.270 -0.035 ;
        RECT 28.270 -0.035 56.565 0.000 ;
      LAYER met2 ;
        RECT 0.500 3.905 74.700 194.395 ;
        RECT 0.500 3.625 54.435 3.905 ;
        RECT 0.500 1.730 54.715 3.625 ;
        RECT 20.775 0.570 54.715 1.730 ;
        RECT 20.775 0.005 34.160 0.570 ;
        RECT 44.720 0.005 54.715 0.570 ;
        RECT 20.775 0.000 34.440 0.005 ;
        RECT 20.925 -0.035 34.440 0.000 ;
        RECT 44.440 0.000 54.715 0.005 ;
        RECT 44.440 -0.035 53.535 0.000 ;
        RECT 54.095 -0.035 54.715 0.000 ;
      LAYER met3 ;
        RECT 0.490 24.215 74.700 197.965 ;
        RECT 24.900 23.265 50.355 24.215 ;
        RECT 24.900 20.585 37.980 23.265 ;
        RECT 24.900 1.695 25.600 20.585 ;
        RECT 37.280 1.695 37.980 20.585 ;
        RECT 49.655 1.695 50.355 23.265 ;
      LAYER met4 ;
        RECT 1.670 173.350 73.330 197.965 ;
        RECT 0.965 93.365 74.035 173.350 ;
        RECT 1.670 67.600 73.330 93.365 ;
        RECT 0.965 66.900 74.035 67.600 ;
        RECT 1.670 61.650 73.330 66.900 ;
        RECT 0.965 61.050 74.035 61.650 ;
        RECT 1.670 55.800 73.330 61.050 ;
        RECT 0.965 55.100 74.035 55.800 ;
        RECT 1.670 49.710 73.330 50.690 ;
        RECT 0.965 44.600 74.035 45.300 ;
        RECT 1.670 39.150 73.330 44.600 ;
        RECT 0.965 38.550 74.035 39.150 ;
        RECT 1.670 34.300 73.330 38.550 ;
        RECT 0.965 33.700 74.035 34.300 ;
        RECT 1.670 29.450 73.330 33.700 ;
        RECT 0.965 28.850 74.035 29.450 ;
        RECT 1.670 23.400 73.330 28.850 ;
        RECT 0.965 22.800 74.035 23.400 ;
        RECT 1.670 17.350 73.330 22.800 ;
        RECT 0.965 16.750 74.035 17.350 ;
        RECT 1.365 12.500 73.635 16.750 ;
        RECT 0.965 11.900 74.035 12.500 ;
        RECT 1.670 6.450 73.330 11.900 ;
        RECT 0.965 5.850 74.035 6.450 ;
        RECT 1.670 0.000 73.330 5.850 ;
      LAYER met5 ;
        RECT 0.000 168.730 75.000 197.965 ;
        RECT 0.000 98.265 8.670 168.730 ;
        RECT 66.270 98.265 75.000 168.730 ;
        RECT 0.000 94.550 75.000 98.265 ;
        RECT 2.870 34.805 72.130 94.550 ;
        RECT 0.000 34.800 75.000 34.805 ;
        RECT 2.870 16.250 72.130 34.800 ;
        RECT 2.565 13.000 72.435 16.250 ;
        RECT 2.870 0.100 72.130 13.000 ;
  END
END sky130_ef_io__vssio_lvc_pad

#--------EOF---------

MACRO sky130_fd_io__signal_5_sym_hv_local_5term
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__signal_5_sym_hv_local_5term ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.955 BY 12.120 ;
  PIN GATE
    ANTENNAGATEAREA 3.400000 ;
    PORT
      LAYER li1 ;
        RECT 3.310 8.925 4.635 9.335 ;
      LAYER mcon ;
        RECT 3.625 9.065 3.795 9.235 ;
        RECT 3.985 9.065 4.155 9.235 ;
      LAYER met1 ;
        RECT 3.515 8.955 4.260 11.795 ;
    END
  END GATE
  PIN NWELLRING
    ANTENNADIFFAREA 24.296999 ;
    PORT
      LAYER nwell ;
        RECT 0.000 10.760 7.955 12.120 ;
        RECT 0.000 1.360 1.360 10.760 ;
        RECT 6.595 1.360 7.955 10.760 ;
        RECT 0.000 0.000 7.955 1.360 ;
      LAYER li1 ;
        RECT 0.330 11.090 7.625 11.790 ;
        RECT 0.330 1.030 1.030 11.090 ;
        RECT 6.925 1.030 7.625 11.090 ;
        RECT 0.330 0.330 7.625 1.030 ;
      LAYER mcon ;
        RECT 1.535 11.355 1.705 11.525 ;
        RECT 1.895 11.355 2.065 11.525 ;
        RECT 2.255 11.355 2.425 11.525 ;
        RECT 2.615 11.355 2.785 11.525 ;
        RECT 2.975 11.355 3.145 11.525 ;
        RECT 4.795 11.355 4.965 11.525 ;
        RECT 5.155 11.355 5.325 11.525 ;
        RECT 5.515 11.355 5.685 11.525 ;
        RECT 5.875 11.355 6.045 11.525 ;
        RECT 6.235 11.355 6.405 11.525 ;
        RECT 0.595 10.005 0.765 10.175 ;
        RECT 0.595 9.645 0.765 9.815 ;
        RECT 0.595 9.285 0.765 9.455 ;
        RECT 0.595 8.925 0.765 9.095 ;
        RECT 0.595 8.565 0.765 8.735 ;
        RECT 0.595 8.205 0.765 8.375 ;
        RECT 0.595 7.845 0.765 8.015 ;
        RECT 0.595 7.485 0.765 7.655 ;
        RECT 0.595 7.125 0.765 7.295 ;
        RECT 0.595 6.765 0.765 6.935 ;
        RECT 0.595 6.405 0.765 6.575 ;
        RECT 0.595 6.045 0.765 6.215 ;
        RECT 0.595 5.685 0.765 5.855 ;
        RECT 0.595 5.325 0.765 5.495 ;
        RECT 0.595 4.965 0.765 5.135 ;
        RECT 0.595 4.605 0.765 4.775 ;
        RECT 0.595 4.245 0.765 4.415 ;
        RECT 0.595 3.885 0.765 4.055 ;
        RECT 0.595 3.525 0.765 3.695 ;
        RECT 0.595 3.165 0.765 3.335 ;
        RECT 0.595 2.805 0.765 2.975 ;
        RECT 0.595 2.445 0.765 2.615 ;
        RECT 0.595 2.085 0.765 2.255 ;
        RECT 0.595 1.725 0.765 1.895 ;
        RECT 0.595 1.365 0.765 1.535 ;
        RECT 7.190 10.005 7.360 10.175 ;
        RECT 7.190 9.645 7.360 9.815 ;
        RECT 7.190 9.285 7.360 9.455 ;
        RECT 7.190 8.925 7.360 9.095 ;
        RECT 7.190 8.565 7.360 8.735 ;
        RECT 7.190 8.205 7.360 8.375 ;
        RECT 7.190 7.845 7.360 8.015 ;
        RECT 7.190 7.485 7.360 7.655 ;
        RECT 7.190 7.125 7.360 7.295 ;
        RECT 7.190 6.765 7.360 6.935 ;
        RECT 7.190 6.405 7.360 6.575 ;
        RECT 7.190 6.045 7.360 6.215 ;
        RECT 7.190 5.685 7.360 5.855 ;
        RECT 7.190 5.325 7.360 5.495 ;
        RECT 7.190 4.965 7.360 5.135 ;
        RECT 7.190 4.605 7.360 4.775 ;
        RECT 7.190 4.245 7.360 4.415 ;
        RECT 7.190 3.885 7.360 4.055 ;
        RECT 7.190 3.525 7.360 3.695 ;
        RECT 7.190 3.165 7.360 3.335 ;
        RECT 7.190 2.805 7.360 2.975 ;
        RECT 7.190 2.445 7.360 2.615 ;
        RECT 7.190 2.085 7.360 2.255 ;
        RECT 7.190 1.725 7.360 1.895 ;
        RECT 7.190 1.365 7.360 1.535 ;
        RECT 5.590 0.540 5.760 0.710 ;
        RECT 5.950 0.540 6.120 0.710 ;
        RECT 6.310 0.540 6.480 0.710 ;
      LAYER met1 ;
        POLYGON 1.040 11.790 1.040 11.080 0.330 11.080 ;
        RECT 1.040 11.090 3.345 11.790 ;
        RECT 4.430 11.090 6.915 11.790 ;
        RECT 1.040 11.080 1.430 11.090 ;
        POLYGON 1.430 11.090 1.440 11.090 1.430 11.080 ;
        POLYGON 6.445 11.090 6.455 11.090 6.455 11.080 ;
        RECT 6.455 11.080 6.915 11.090 ;
        POLYGON 6.915 11.790 7.625 11.080 6.915 11.080 ;
        RECT 0.330 0.345 1.030 11.080 ;
        POLYGON 1.030 11.080 1.430 11.080 1.030 10.680 ;
        POLYGON 6.455 11.080 6.855 11.080 6.855 10.680 ;
        RECT 6.855 10.680 7.625 11.080 ;
        POLYGON 6.855 10.680 6.915 10.680 6.915 10.620 ;
        RECT 6.915 10.620 7.625 10.680 ;
        POLYGON 6.915 10.620 6.925 10.620 6.925 10.610 ;
        POLYGON 6.925 1.510 6.925 1.030 6.445 1.030 ;
        RECT 6.925 1.040 7.625 10.620 ;
        RECT 6.925 1.030 6.930 1.040 ;
        RECT 5.350 0.345 6.930 1.030 ;
        POLYGON 6.930 1.040 7.625 1.040 6.930 0.345 ;
        RECT 0.330 0.330 1.015 0.345 ;
        RECT 5.350 0.330 6.915 0.345 ;
        POLYGON 6.915 0.345 6.930 0.345 6.915 0.330 ;
    END
  END NWELLRING
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 2.965 3.360 3.505 8.755 ;
      LAYER mcon ;
        RECT 3.105 7.745 3.275 7.915 ;
        RECT 3.105 7.385 3.275 7.555 ;
        RECT 3.105 7.025 3.275 7.195 ;
        RECT 3.105 6.665 3.275 6.835 ;
        RECT 3.105 6.305 3.275 6.475 ;
        RECT 3.105 5.945 3.275 6.115 ;
        RECT 3.105 5.585 3.275 5.755 ;
        RECT 3.105 5.225 3.275 5.395 ;
        RECT 3.105 4.865 3.275 5.035 ;
        RECT 3.105 4.505 3.275 4.675 ;
        RECT 3.105 4.145 3.275 4.315 ;
        RECT 3.105 3.785 3.275 3.955 ;
      LAYER met1 ;
        RECT 2.860 0.330 3.860 8.545 ;
    END
  END VGND
  PIN NBODY
    ANTENNADIFFAREA 13.550600 ;
    PORT
      LAYER pwell ;
        RECT 1.660 1.660 6.295 10.460 ;
      LAYER li1 ;
        RECT 1.790 9.620 6.165 10.330 ;
        RECT 1.790 2.490 2.490 9.620 ;
        RECT 5.465 2.490 6.165 9.620 ;
        RECT 1.790 1.790 6.165 2.490 ;
      LAYER mcon ;
        RECT 2.270 9.845 2.440 10.015 ;
        RECT 2.630 9.845 2.800 10.015 ;
        RECT 2.990 9.845 3.160 10.015 ;
        RECT 4.640 9.845 4.810 10.015 ;
        RECT 5.000 9.845 5.170 10.015 ;
        RECT 5.360 9.845 5.530 10.015 ;
        RECT 1.975 8.845 2.145 9.015 ;
        RECT 1.975 8.485 2.145 8.655 ;
        RECT 1.975 8.125 2.145 8.295 ;
        RECT 1.975 7.765 2.145 7.935 ;
        RECT 1.975 7.405 2.145 7.575 ;
        RECT 1.975 7.045 2.145 7.215 ;
        RECT 1.975 6.685 2.145 6.855 ;
        RECT 1.975 6.325 2.145 6.495 ;
        RECT 1.975 5.965 2.145 6.135 ;
        RECT 1.975 5.605 2.145 5.775 ;
        RECT 1.975 5.245 2.145 5.415 ;
        RECT 1.975 4.885 2.145 5.055 ;
        RECT 1.975 4.525 2.145 4.695 ;
        RECT 1.975 4.165 2.145 4.335 ;
        RECT 1.975 3.805 2.145 3.975 ;
        RECT 1.975 3.445 2.145 3.615 ;
        RECT 1.975 3.085 2.145 3.255 ;
        RECT 1.975 2.725 2.145 2.895 ;
        RECT 1.975 2.365 2.145 2.535 ;
        RECT 5.730 8.845 5.900 9.015 ;
        RECT 5.730 8.485 5.900 8.655 ;
        RECT 5.730 8.125 5.900 8.295 ;
        RECT 5.730 7.765 5.900 7.935 ;
        RECT 5.730 7.405 5.900 7.575 ;
        RECT 5.730 7.045 5.900 7.215 ;
        RECT 5.730 6.685 5.900 6.855 ;
        RECT 5.730 6.325 5.900 6.495 ;
        RECT 5.730 5.965 5.900 6.135 ;
        RECT 5.730 5.605 5.900 5.775 ;
        RECT 5.730 5.245 5.900 5.415 ;
        RECT 5.730 4.885 5.900 5.055 ;
        RECT 5.730 4.525 5.900 4.695 ;
        RECT 5.730 4.165 5.900 4.335 ;
        RECT 5.730 3.805 5.900 3.975 ;
        RECT 5.730 3.445 5.900 3.615 ;
        RECT 5.730 3.085 5.900 3.255 ;
        RECT 5.730 2.725 5.900 2.895 ;
        RECT 5.730 2.365 5.900 2.535 ;
        RECT 1.975 2.005 2.145 2.175 ;
        RECT 5.730 2.005 5.900 2.175 ;
      LAYER met1 ;
        POLYGON 2.120 10.330 2.120 10.000 1.790 10.000 ;
        RECT 2.120 10.000 3.345 10.330 ;
        RECT 1.790 9.505 3.345 10.000 ;
        RECT 4.430 10.000 5.835 10.330 ;
        POLYGON 5.835 10.330 6.165 10.000 5.835 10.000 ;
        RECT 4.430 9.505 6.165 10.000 ;
        RECT 1.790 0.345 2.680 9.505 ;
        POLYGON 2.680 9.505 3.055 9.505 2.680 9.130 ;
        POLYGON 5.060 9.505 5.435 9.505 5.435 9.130 ;
        RECT 5.435 9.130 6.165 9.505 ;
        POLYGON 5.435 9.130 5.465 9.130 5.465 9.100 ;
        RECT 5.465 1.790 6.165 9.130 ;
        RECT 1.790 0.330 2.665 0.345 ;
    END
  END NBODY
  PIN IN
    ANTENNADIFFAREA 3.807000 ;
    PORT
      LAYER li1 ;
        RECT 4.440 3.360 4.980 8.755 ;
      LAYER mcon ;
        RECT 4.575 7.745 4.745 7.915 ;
        RECT 4.575 7.385 4.745 7.555 ;
        RECT 4.575 7.025 4.745 7.195 ;
        RECT 4.575 6.665 4.745 6.835 ;
        RECT 4.575 6.305 4.745 6.475 ;
        RECT 4.575 5.945 4.745 6.115 ;
        RECT 4.575 5.585 4.745 5.755 ;
        RECT 4.575 5.225 4.745 5.395 ;
        RECT 4.575 4.865 4.745 5.035 ;
        RECT 4.575 4.505 4.745 4.675 ;
        RECT 4.575 4.145 4.745 4.315 ;
        RECT 4.575 3.785 4.745 3.955 ;
      LAYER met1 ;
        RECT 4.155 0.330 5.155 8.760 ;
    END
  END IN
  OBS
      LAYER met1 ;
        RECT 1.015 0.330 1.030 0.345 ;
        RECT 2.665 0.330 2.680 0.345 ;
  END
END sky130_fd_io__signal_5_sym_hv_local_5term

#--------EOF---------


END LIBRARY
